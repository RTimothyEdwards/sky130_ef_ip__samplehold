magic
tech sky130A
magscale 1 2
timestamp 1652202333
<< locali >>
rect 392 8914 616 9238
rect 940 9208 2054 9238
rect 940 8946 1166 9208
rect 2008 8946 2054 9208
rect 940 8914 2054 8946
rect 392 8734 426 8914
rect 2020 8732 2054 8914
rect 722 8622 830 8646
rect 722 8262 744 8622
rect 814 8262 830 8622
rect 722 8214 830 8262
rect 1692 6610 1778 6648
rect 1428 6600 1778 6610
rect 1428 6536 1440 6600
rect 1764 6536 1778 6600
rect 1428 6524 1778 6536
<< viali >>
rect 1166 8946 2008 9208
rect 744 8262 814 8622
rect 1440 6536 1764 6600
<< metal1 >>
rect 11011 11170 11403 11182
rect 11011 10890 11023 11170
rect 11389 10890 11403 11170
rect 11011 10153 11403 10890
rect 0 9612 1070 9952
rect 0 9040 200 9101
rect 0 8950 815 9040
rect 0 8901 200 8950
rect 743 8632 815 8950
rect 1013 8655 1070 9612
rect 1118 9208 2060 9238
rect 1118 8946 1166 9208
rect 2008 8946 2060 9208
rect 1118 8914 2060 8946
rect 1912 8702 1986 8914
rect 2014 8738 2060 8914
rect 2014 8702 2020 8738
rect 2054 8702 2060 8738
rect 732 8622 826 8632
rect 732 8262 744 8622
rect 814 8262 826 8622
rect 732 8246 826 8262
rect 386 6474 432 6652
rect 460 6474 534 6652
rect 0 6462 1040 6474
rect 0 6166 814 6462
rect 1026 6166 1040 6462
rect 0 6152 1040 6166
rect 1098 6082 1172 6700
rect 1200 6082 1246 6646
rect 1274 6082 1348 6700
rect 1428 6600 1778 6610
rect 1428 6536 1440 6600
rect 1764 6536 1778 6600
rect 1428 6524 1778 6536
rect 1912 6476 1986 6640
rect 2014 6476 2060 6640
rect 1406 6464 2060 6476
rect 1406 6168 1422 6464
rect 1616 6168 2060 6464
rect 1406 6152 2060 6168
rect 11011 6327 11403 9266
rect 1098 6015 1348 6082
rect 0 5284 2515 6015
rect 3391 5284 3424 6015
rect 11011 5969 11029 6327
rect 11387 5969 11403 6327
rect 11011 5949 11403 5969
rect 10725 5488 12368 5842
rect 11011 5340 11403 5360
rect 0 4986 3717 5186
rect 11011 4982 11028 5340
rect 11386 4982 11403 5340
rect 0 4641 1888 4841
rect 2381 4641 3717 4841
rect 11011 4451 11403 4982
rect 2404 2443 2515 2719
rect 3391 2443 3517 2719
rect 2924 1925 3657 2298
rect 11011 2289 11403 4050
rect 2416 1647 2693 1847
rect 2493 1595 2693 1647
rect 2493 1427 2693 1436
rect 2924 1287 3506 1925
rect 2924 941 2942 1287
rect 2402 726 2942 941
rect 3484 726 3506 1287
rect 2402 706 3506 726
rect 11011 627 11403 660
rect 11546 4996 12150 5196
rect 11546 281 11746 4996
rect 11875 4651 12150 4851
rect 11875 483 11987 4651
rect 19130 4570 19469 4770
rect 11875 370 11885 483
rect 12206 370 12216 483
rect 2478 248 3021 281
rect 2478 -80 2519 248
rect 2985 -80 3021 248
rect 2478 -114 3021 -80
rect 11278 248 11821 281
rect 11278 -80 11319 248
rect 11785 -80 11821 248
rect 11278 -114 11821 -80
<< via1 >>
rect 11023 10890 11389 11170
rect 11011 9266 11403 10153
rect 814 6166 1026 6462
rect 1440 6536 1764 6600
rect 1422 6168 1616 6464
rect 2515 5284 3391 6015
rect 11029 5969 11387 6327
rect 11028 4982 11386 5340
rect 1888 4641 2381 4841
rect 11011 4050 11403 4451
rect 2515 2443 3391 2719
rect 2493 1436 2693 1595
rect 872 718 1589 929
rect 2942 726 3484 1287
rect 11011 660 11403 2289
rect 11885 370 12206 483
rect 2519 -80 2985 248
rect 11319 -80 11785 248
<< metal2 >>
rect 11011 11170 11403 11182
rect 2515 10932 3391 11027
rect 2515 10710 3685 10932
rect 10732 10756 10958 10932
rect 11011 10890 11023 11170
rect 11389 10890 11403 11170
rect 11011 10836 11403 10890
rect 11477 10756 12149 10942
rect 10732 10710 12149 10756
rect 1428 6600 1778 6610
rect 1428 6536 1440 6600
rect 1764 6536 1778 6600
rect 1428 6524 1778 6536
rect 798 6464 1630 6474
rect 798 6462 1422 6464
rect 798 6166 814 6462
rect 1026 6168 1422 6462
rect 1616 6168 1630 6464
rect 1026 6166 1630 6168
rect 798 6152 1630 6166
rect 1692 3414 1778 6524
rect 2515 6015 3391 10710
rect 10835 10479 11721 10710
rect 11011 10153 11403 10231
rect 11011 6327 11403 9266
rect 11011 5969 11029 6327
rect 11387 5969 11403 6327
rect 3391 5573 3685 5842
rect 1871 4641 1888 4841
rect 2381 4641 2394 4841
rect 856 929 1605 940
rect 856 718 872 929
rect 1589 718 1605 929
rect 856 706 1605 718
rect 2300 464 2394 4641
rect 2515 2719 3391 5284
rect 11011 5340 11403 5969
rect 11011 4982 11028 5340
rect 11386 4982 11403 5340
rect 2515 2403 3391 2443
rect 10573 1595 10732 4882
rect 11011 4451 11403 4982
rect 10976 4050 11011 4451
rect 11403 4050 12119 4451
rect 2484 1436 2493 1595
rect 2693 1436 10732 1595
rect 10952 2289 12119 2326
rect 2924 1287 3506 1305
rect 2924 726 2942 1287
rect 3484 803 3506 1287
rect 10952 803 11011 2289
rect 3484 726 11011 803
rect 2924 660 11011 726
rect 11403 1934 12119 2289
rect 11403 803 11921 1934
rect 11403 660 19235 803
rect 2924 578 19235 660
rect 11875 464 11885 483
rect 2300 370 11885 464
rect 12206 370 12216 483
rect 2478 248 3021 281
rect 2478 -80 2519 248
rect 2985 -80 3021 248
rect 2478 -114 3021 -80
rect 11278 248 11821 281
rect 11278 -80 11319 248
rect 11785 -80 11821 248
rect 11278 -114 11821 -80
<< via2 >>
rect 11023 10890 11389 11170
rect 357 1087 508 2307
rect 872 718 1589 929
rect 2519 -80 2985 248
rect 11319 -80 11785 248
<< metal3 >>
rect 11011 11170 11403 11182
rect 11011 10890 11023 11170
rect 11389 10890 11403 11170
rect 11011 10879 11403 10890
rect 337 2307 522 2321
rect 337 1087 357 2307
rect 508 1087 522 2307
rect 337 191 522 1087
rect 856 929 1605 940
rect 856 718 872 929
rect 1589 718 1605 929
rect 856 706 1605 718
rect 2478 248 3021 281
rect 2478 191 2519 248
rect 337 6 2519 191
rect 2478 -80 2519 6
rect 2985 -80 3021 248
rect 2478 -114 3021 -80
rect 11278 248 11821 281
rect 11278 -80 11319 248
rect 11785 -80 11821 248
rect 11278 -114 11821 -80
<< via3 >>
rect 11023 10890 11389 11170
rect 872 718 1589 929
rect 2519 -80 2985 248
rect 11319 -80 11785 248
<< metal4 >>
rect 0 11182 1039 11183
rect 0 10817 2236 11182
rect 0 10191 1606 10817
rect 857 929 1606 10191
rect 857 718 872 929
rect 1589 718 1606 929
rect 857 637 1606 718
rect 2478 248 3021 281
rect 2478 -80 2519 248
rect 2985 -80 3021 248
rect 2478 -114 3021 -80
rect 11278 248 11821 281
rect 11278 -80 11319 248
rect 11785 -80 11821 248
rect 11278 -114 11821 -80
<< via4 >>
rect 2519 -80 2985 248
rect 11319 -80 11785 248
<< metal5 >>
rect 2478 248 3021 281
rect 2478 -80 2519 248
rect 2985 -80 3021 248
rect 2478 -114 3021 -80
rect 11278 248 11871 281
rect 11278 -80 11319 248
rect 11785 -80 11871 248
rect 11278 -114 11871 -80
use hold_cap_array  hold_cap_array_0
timestamp 1652200182
transform 1 0 218 0 1 26439
box 1997 -26553 19047 -15257
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_0 paramcells
timestamp 1652200182
transform 1 0 778 0 1 9076
box -198 -198 198 198
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1650294714
transform 0 1 409 -1 0 8738
box -66 -43 2178 1671
use balanced_switch  x1
timestamp 1652200182
transform -1 0 2730 0 1 2811
box 301 -2311 2543 1830
use follower_amp  x2
timestamp 1652202333
transform 1 0 8047 0 1 4397
box -4547 -3901 2817 6641
use follower_amp  x3
timestamp 1652202333
transform 1 0 16511 0 1 4407
box -4547 -3901 2817 6641
<< labels >>
flabel metal1 0 5284 200 6015 0 FreeSans 320 0 0 0 vdd
port 2 nsew
flabel metal1 0 8901 200 9101 0 FreeSans 256 0 0 0 hold
port 3 nsew
flabel metal1 0 9612 804 9952 0 FreeSans 1600 0 0 0 dvdd
port 6 nsew
flabel metal1 0 6152 788 6474 0 FreeSans 1600 0 0 0 dvss
port 7 nsew
flabel metal4 0 10191 1039 11183 0 FreeSans 1600 0 0 0 vss
port 5 nsew
flabel metal1 19269 4570 19469 4770 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 0 4986 200 5186 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal1 0 4641 200 4841 0 FreeSans 320 0 0 0 ena
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 19469 11297
<< end >>
