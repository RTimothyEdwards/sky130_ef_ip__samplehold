magic
tech sky130A
magscale 1 2
timestamp 1651944383
<< error_p >>
rect -111 10234 -91 10400
rect 209 10234 229 10400
rect -111 8934 -91 9266
rect 209 8934 229 9266
rect -111 7634 -91 7966
rect 209 7634 229 7966
rect -111 6334 -91 6666
rect 209 6334 229 6666
rect -111 5034 -91 5366
rect 209 5034 229 5366
rect -111 3734 -91 4066
rect 209 3734 229 4066
rect -111 2434 -91 2766
rect 209 2434 229 2766
rect -111 1134 -91 1466
rect 209 1134 229 1466
rect -111 -166 -91 166
rect 209 -166 229 166
rect -111 -1466 -91 -1134
rect 209 -1466 229 -1134
rect -111 -2766 -91 -2434
rect 209 -2766 229 -2434
rect -111 -4066 -91 -3734
rect 209 -4066 229 -3734
rect -111 -5366 -91 -5034
rect 209 -5366 229 -5034
rect -111 -6666 -91 -6334
rect 209 -6666 229 -6334
rect -111 -7966 -91 -7634
rect 209 -7966 229 -7634
rect -111 -9266 -91 -8934
rect 209 -9266 229 -8934
rect -111 -10400 -91 -10234
rect 209 -10400 229 -10234
rect 233 -10400 529 10400
rect 553 9371 849 10351
rect 553 9149 873 9371
rect 553 8829 873 9051
rect 553 8071 849 8829
rect 553 7849 873 8071
rect 553 7529 873 7751
rect 553 6771 849 7529
rect 553 6549 873 6771
rect 553 6229 873 6451
rect 553 5471 849 6229
rect 553 5249 873 5471
rect 553 4929 873 5151
rect 553 4171 849 4929
rect 553 3949 873 4171
rect 553 3629 873 3851
rect 553 2871 849 3629
rect 553 2649 873 2871
rect 553 2329 873 2551
rect 553 1571 849 2329
rect 553 1349 873 1571
rect 553 1029 873 1251
rect 553 271 849 1029
rect 553 49 873 271
rect 553 -271 873 -49
rect 553 -1029 849 -271
rect 553 -1251 873 -1029
rect 553 -1571 873 -1349
rect 553 -2329 849 -1571
rect 553 -2551 873 -2329
rect 553 -2871 873 -2649
rect 553 -3629 849 -2871
rect 553 -3851 873 -3629
rect 553 -4171 873 -3949
rect 553 -4929 849 -4171
rect 553 -5151 873 -4929
rect 553 -5471 873 -5249
rect 553 -6229 849 -5471
rect 553 -6451 873 -6229
rect 553 -6771 873 -6549
rect 553 -7529 849 -6771
rect 553 -7751 873 -7529
rect 553 -8071 873 -7849
rect 553 -8829 849 -8071
rect 553 -9051 873 -8829
rect 553 -9371 873 -9149
rect 553 -10351 849 -9371
<< metal4 >>
rect -851 10309 851 10350
rect -851 9191 595 10309
rect 831 9191 851 10309
rect -851 9150 851 9191
rect -851 9009 851 9050
rect -851 7891 595 9009
rect 831 7891 851 9009
rect -851 7850 851 7891
rect -851 7709 851 7750
rect -851 6591 595 7709
rect 831 6591 851 7709
rect -851 6550 851 6591
rect -851 6409 851 6450
rect -851 5291 595 6409
rect 831 5291 851 6409
rect -851 5250 851 5291
rect -851 5109 851 5150
rect -851 3991 595 5109
rect 831 3991 851 5109
rect -851 3950 851 3991
rect -851 3809 851 3850
rect -851 2691 595 3809
rect 831 2691 851 3809
rect -851 2650 851 2691
rect -851 2509 851 2550
rect -851 1391 595 2509
rect 831 1391 851 2509
rect -851 1350 851 1391
rect -851 1209 851 1250
rect -851 91 595 1209
rect 831 91 851 1209
rect -851 50 851 91
rect -851 -91 851 -50
rect -851 -1209 595 -91
rect 831 -1209 851 -91
rect -851 -1250 851 -1209
rect -851 -1391 851 -1350
rect -851 -2509 595 -1391
rect 831 -2509 851 -1391
rect -851 -2550 851 -2509
rect -851 -2691 851 -2650
rect -851 -3809 595 -2691
rect 831 -3809 851 -2691
rect -851 -3850 851 -3809
rect -851 -3991 851 -3950
rect -851 -5109 595 -3991
rect 831 -5109 851 -3991
rect -851 -5150 851 -5109
rect -851 -5291 851 -5250
rect -851 -6409 595 -5291
rect 831 -6409 851 -5291
rect -851 -6450 851 -6409
rect -851 -6591 851 -6550
rect -851 -7709 595 -6591
rect 831 -7709 851 -6591
rect -851 -7750 851 -7709
rect -851 -7891 851 -7850
rect -851 -9009 595 -7891
rect 831 -9009 851 -7891
rect -851 -9050 851 -9009
rect -851 -9191 851 -9150
rect -851 -10309 595 -9191
rect 831 -10309 851 -9191
rect -851 -10350 851 -10309
<< via4 >>
rect 595 9191 831 10309
rect 595 7891 831 9009
rect 595 6591 831 7709
rect 595 5291 831 6409
rect 595 3991 831 5109
rect 595 2691 831 3809
rect 595 1391 831 2509
rect 595 91 831 1209
rect 595 -1209 831 -91
rect 595 -2509 831 -1391
rect 595 -3809 831 -2691
rect 595 -5109 831 -3991
rect 595 -6409 831 -5291
rect 595 -7709 831 -6591
rect 595 -9009 831 -7891
rect 595 -10309 831 -9191
<< mimcap2 >>
rect -751 10210 249 10250
rect -751 9290 -711 10210
rect 209 9290 249 10210
rect -751 9250 249 9290
rect -751 8910 249 8950
rect -751 7990 -711 8910
rect 209 7990 249 8910
rect -751 7950 249 7990
rect -751 7610 249 7650
rect -751 6690 -711 7610
rect 209 6690 249 7610
rect -751 6650 249 6690
rect -751 6310 249 6350
rect -751 5390 -711 6310
rect 209 5390 249 6310
rect -751 5350 249 5390
rect -751 5010 249 5050
rect -751 4090 -711 5010
rect 209 4090 249 5010
rect -751 4050 249 4090
rect -751 3710 249 3750
rect -751 2790 -711 3710
rect 209 2790 249 3710
rect -751 2750 249 2790
rect -751 2410 249 2450
rect -751 1490 -711 2410
rect 209 1490 249 2410
rect -751 1450 249 1490
rect -751 1110 249 1150
rect -751 190 -711 1110
rect 209 190 249 1110
rect -751 150 249 190
rect -751 -190 249 -150
rect -751 -1110 -711 -190
rect 209 -1110 249 -190
rect -751 -1150 249 -1110
rect -751 -1490 249 -1450
rect -751 -2410 -711 -1490
rect 209 -2410 249 -1490
rect -751 -2450 249 -2410
rect -751 -2790 249 -2750
rect -751 -3710 -711 -2790
rect 209 -3710 249 -2790
rect -751 -3750 249 -3710
rect -751 -4090 249 -4050
rect -751 -5010 -711 -4090
rect 209 -5010 249 -4090
rect -751 -5050 249 -5010
rect -751 -5390 249 -5350
rect -751 -6310 -711 -5390
rect 209 -6310 249 -5390
rect -751 -6350 249 -6310
rect -751 -6690 249 -6650
rect -751 -7610 -711 -6690
rect 209 -7610 249 -6690
rect -751 -7650 249 -7610
rect -751 -7990 249 -7950
rect -751 -8910 -711 -7990
rect 209 -8910 249 -7990
rect -751 -8950 249 -8910
rect -751 -9290 249 -9250
rect -751 -10210 -711 -9290
rect 209 -10210 249 -9290
rect -751 -10250 249 -10210
<< mimcap2contact >>
rect -711 9290 209 10210
rect -711 7990 209 8910
rect -711 6690 209 7610
rect -711 5390 209 6310
rect -711 4090 209 5010
rect -711 2790 209 3710
rect -711 1490 209 2410
rect -711 190 209 1110
rect -711 -1110 209 -190
rect -711 -2410 209 -1490
rect -711 -3710 209 -2790
rect -711 -5010 209 -4090
rect -711 -6310 209 -5390
rect -711 -7610 209 -6690
rect -711 -8910 209 -7990
rect -711 -10210 209 -9290
<< metal5 >>
rect -411 10234 -91 10400
rect 209 10234 529 10400
rect -735 10210 529 10234
rect -735 9290 -711 10210
rect 209 9290 529 10210
rect -735 9266 529 9290
rect -411 8934 -91 9266
rect 209 8934 529 9266
rect 553 10309 873 10351
rect 553 9191 595 10309
rect 831 9191 873 10309
rect 553 9149 873 9191
rect -735 8910 529 8934
rect -735 7990 -711 8910
rect 209 7990 529 8910
rect -735 7966 529 7990
rect -411 7634 -91 7966
rect 209 7634 529 7966
rect 553 9009 873 9051
rect 553 7891 595 9009
rect 831 7891 873 9009
rect 553 7849 873 7891
rect -735 7610 529 7634
rect -735 6690 -711 7610
rect 209 6690 529 7610
rect -735 6666 529 6690
rect -411 6334 -91 6666
rect 209 6334 529 6666
rect 553 7709 873 7751
rect 553 6591 595 7709
rect 831 6591 873 7709
rect 553 6549 873 6591
rect -735 6310 529 6334
rect -735 5390 -711 6310
rect 209 5390 529 6310
rect -735 5366 529 5390
rect -411 5034 -91 5366
rect 209 5034 529 5366
rect 553 6409 873 6451
rect 553 5291 595 6409
rect 831 5291 873 6409
rect 553 5249 873 5291
rect -735 5010 529 5034
rect -735 4090 -711 5010
rect 209 4090 529 5010
rect -735 4066 529 4090
rect -411 3734 -91 4066
rect 209 3734 529 4066
rect 553 5109 873 5151
rect 553 3991 595 5109
rect 831 3991 873 5109
rect 553 3949 873 3991
rect -735 3710 529 3734
rect -735 2790 -711 3710
rect 209 2790 529 3710
rect -735 2766 529 2790
rect -411 2434 -91 2766
rect 209 2434 529 2766
rect 553 3809 873 3851
rect 553 2691 595 3809
rect 831 2691 873 3809
rect 553 2649 873 2691
rect -735 2410 529 2434
rect -735 1490 -711 2410
rect 209 1490 529 2410
rect -735 1466 529 1490
rect -411 1134 -91 1466
rect 209 1134 529 1466
rect 553 2509 873 2551
rect 553 1391 595 2509
rect 831 1391 873 2509
rect 553 1349 873 1391
rect -735 1110 529 1134
rect -735 190 -711 1110
rect 209 190 529 1110
rect -735 166 529 190
rect -411 -166 -91 166
rect 209 -166 529 166
rect 553 1209 873 1251
rect 553 91 595 1209
rect 831 91 873 1209
rect 553 49 873 91
rect -735 -190 529 -166
rect -735 -1110 -711 -190
rect 209 -1110 529 -190
rect -735 -1134 529 -1110
rect -411 -1466 -91 -1134
rect 209 -1466 529 -1134
rect 553 -91 873 -49
rect 553 -1209 595 -91
rect 831 -1209 873 -91
rect 553 -1251 873 -1209
rect -735 -1490 529 -1466
rect -735 -2410 -711 -1490
rect 209 -2410 529 -1490
rect -735 -2434 529 -2410
rect -411 -2766 -91 -2434
rect 209 -2766 529 -2434
rect 553 -1391 873 -1349
rect 553 -2509 595 -1391
rect 831 -2509 873 -1391
rect 553 -2551 873 -2509
rect -735 -2790 529 -2766
rect -735 -3710 -711 -2790
rect 209 -3710 529 -2790
rect -735 -3734 529 -3710
rect -411 -4066 -91 -3734
rect 209 -4066 529 -3734
rect 553 -2691 873 -2649
rect 553 -3809 595 -2691
rect 831 -3809 873 -2691
rect 553 -3851 873 -3809
rect -735 -4090 529 -4066
rect -735 -5010 -711 -4090
rect 209 -5010 529 -4090
rect -735 -5034 529 -5010
rect -411 -5366 -91 -5034
rect 209 -5366 529 -5034
rect 553 -3991 873 -3949
rect 553 -5109 595 -3991
rect 831 -5109 873 -3991
rect 553 -5151 873 -5109
rect -735 -5390 529 -5366
rect -735 -6310 -711 -5390
rect 209 -6310 529 -5390
rect -735 -6334 529 -6310
rect -411 -6666 -91 -6334
rect 209 -6666 529 -6334
rect 553 -5291 873 -5249
rect 553 -6409 595 -5291
rect 831 -6409 873 -5291
rect 553 -6451 873 -6409
rect -735 -6690 529 -6666
rect -735 -7610 -711 -6690
rect 209 -7610 529 -6690
rect -735 -7634 529 -7610
rect -411 -7966 -91 -7634
rect 209 -7966 529 -7634
rect 553 -6591 873 -6549
rect 553 -7709 595 -6591
rect 831 -7709 873 -6591
rect 553 -7751 873 -7709
rect -735 -7990 529 -7966
rect -735 -8910 -711 -7990
rect 209 -8910 529 -7990
rect -735 -8934 529 -8910
rect -411 -9266 -91 -8934
rect 209 -9266 529 -8934
rect 553 -7891 873 -7849
rect 553 -9009 595 -7891
rect 831 -9009 873 -7891
rect 553 -9051 873 -9009
rect -735 -9290 529 -9266
rect -735 -10210 -711 -9290
rect 209 -10210 529 -9290
rect -735 -10234 529 -10210
rect -411 -10400 -91 -10234
rect 209 -10400 529 -10234
rect 553 -9191 873 -9149
rect 553 -10309 595 -9191
rect 831 -10309 873 -9191
rect 553 -10351 873 -10309
<< properties >>
string FIXED_BBOX -851 9150 349 10350
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 1 ny 16 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
