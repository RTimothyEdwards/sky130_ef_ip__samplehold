magic
tech sky130A
magscale 1 2
timestamp 1717690002
<< nwell >>
rect -2441 -2359 2441 2359
<< mvpmos >>
rect -2183 1862 -2083 2062
rect -2025 1862 -1925 2062
rect -1867 1862 -1767 2062
rect -1709 1862 -1609 2062
rect -1551 1862 -1451 2062
rect -1393 1862 -1293 2062
rect -1235 1862 -1135 2062
rect -1077 1862 -977 2062
rect -919 1862 -819 2062
rect -761 1862 -661 2062
rect -603 1862 -503 2062
rect -445 1862 -345 2062
rect -287 1862 -187 2062
rect -129 1862 -29 2062
rect 29 1862 129 2062
rect 187 1862 287 2062
rect 345 1862 445 2062
rect 503 1862 603 2062
rect 661 1862 761 2062
rect 819 1862 919 2062
rect 977 1862 1077 2062
rect 1135 1862 1235 2062
rect 1293 1862 1393 2062
rect 1451 1862 1551 2062
rect 1609 1862 1709 2062
rect 1767 1862 1867 2062
rect 1925 1862 2025 2062
rect 2083 1862 2183 2062
rect -2183 1426 -2083 1626
rect -2025 1426 -1925 1626
rect -1867 1426 -1767 1626
rect -1709 1426 -1609 1626
rect -1551 1426 -1451 1626
rect -1393 1426 -1293 1626
rect -1235 1426 -1135 1626
rect -1077 1426 -977 1626
rect -919 1426 -819 1626
rect -761 1426 -661 1626
rect -603 1426 -503 1626
rect -445 1426 -345 1626
rect -287 1426 -187 1626
rect -129 1426 -29 1626
rect 29 1426 129 1626
rect 187 1426 287 1626
rect 345 1426 445 1626
rect 503 1426 603 1626
rect 661 1426 761 1626
rect 819 1426 919 1626
rect 977 1426 1077 1626
rect 1135 1426 1235 1626
rect 1293 1426 1393 1626
rect 1451 1426 1551 1626
rect 1609 1426 1709 1626
rect 1767 1426 1867 1626
rect 1925 1426 2025 1626
rect 2083 1426 2183 1626
rect -2183 990 -2083 1190
rect -2025 990 -1925 1190
rect -1867 990 -1767 1190
rect -1709 990 -1609 1190
rect -1551 990 -1451 1190
rect -1393 990 -1293 1190
rect -1235 990 -1135 1190
rect -1077 990 -977 1190
rect -919 990 -819 1190
rect -761 990 -661 1190
rect -603 990 -503 1190
rect -445 990 -345 1190
rect -287 990 -187 1190
rect -129 990 -29 1190
rect 29 990 129 1190
rect 187 990 287 1190
rect 345 990 445 1190
rect 503 990 603 1190
rect 661 990 761 1190
rect 819 990 919 1190
rect 977 990 1077 1190
rect 1135 990 1235 1190
rect 1293 990 1393 1190
rect 1451 990 1551 1190
rect 1609 990 1709 1190
rect 1767 990 1867 1190
rect 1925 990 2025 1190
rect 2083 990 2183 1190
rect -2183 554 -2083 754
rect -2025 554 -1925 754
rect -1867 554 -1767 754
rect -1709 554 -1609 754
rect -1551 554 -1451 754
rect -1393 554 -1293 754
rect -1235 554 -1135 754
rect -1077 554 -977 754
rect -919 554 -819 754
rect -761 554 -661 754
rect -603 554 -503 754
rect -445 554 -345 754
rect -287 554 -187 754
rect -129 554 -29 754
rect 29 554 129 754
rect 187 554 287 754
rect 345 554 445 754
rect 503 554 603 754
rect 661 554 761 754
rect 819 554 919 754
rect 977 554 1077 754
rect 1135 554 1235 754
rect 1293 554 1393 754
rect 1451 554 1551 754
rect 1609 554 1709 754
rect 1767 554 1867 754
rect 1925 554 2025 754
rect 2083 554 2183 754
rect -2183 118 -2083 318
rect -2025 118 -1925 318
rect -1867 118 -1767 318
rect -1709 118 -1609 318
rect -1551 118 -1451 318
rect -1393 118 -1293 318
rect -1235 118 -1135 318
rect -1077 118 -977 318
rect -919 118 -819 318
rect -761 118 -661 318
rect -603 118 -503 318
rect -445 118 -345 318
rect -287 118 -187 318
rect -129 118 -29 318
rect 29 118 129 318
rect 187 118 287 318
rect 345 118 445 318
rect 503 118 603 318
rect 661 118 761 318
rect 819 118 919 318
rect 977 118 1077 318
rect 1135 118 1235 318
rect 1293 118 1393 318
rect 1451 118 1551 318
rect 1609 118 1709 318
rect 1767 118 1867 318
rect 1925 118 2025 318
rect 2083 118 2183 318
rect -2183 -318 -2083 -118
rect -2025 -318 -1925 -118
rect -1867 -318 -1767 -118
rect -1709 -318 -1609 -118
rect -1551 -318 -1451 -118
rect -1393 -318 -1293 -118
rect -1235 -318 -1135 -118
rect -1077 -318 -977 -118
rect -919 -318 -819 -118
rect -761 -318 -661 -118
rect -603 -318 -503 -118
rect -445 -318 -345 -118
rect -287 -318 -187 -118
rect -129 -318 -29 -118
rect 29 -318 129 -118
rect 187 -318 287 -118
rect 345 -318 445 -118
rect 503 -318 603 -118
rect 661 -318 761 -118
rect 819 -318 919 -118
rect 977 -318 1077 -118
rect 1135 -318 1235 -118
rect 1293 -318 1393 -118
rect 1451 -318 1551 -118
rect 1609 -318 1709 -118
rect 1767 -318 1867 -118
rect 1925 -318 2025 -118
rect 2083 -318 2183 -118
rect -2183 -754 -2083 -554
rect -2025 -754 -1925 -554
rect -1867 -754 -1767 -554
rect -1709 -754 -1609 -554
rect -1551 -754 -1451 -554
rect -1393 -754 -1293 -554
rect -1235 -754 -1135 -554
rect -1077 -754 -977 -554
rect -919 -754 -819 -554
rect -761 -754 -661 -554
rect -603 -754 -503 -554
rect -445 -754 -345 -554
rect -287 -754 -187 -554
rect -129 -754 -29 -554
rect 29 -754 129 -554
rect 187 -754 287 -554
rect 345 -754 445 -554
rect 503 -754 603 -554
rect 661 -754 761 -554
rect 819 -754 919 -554
rect 977 -754 1077 -554
rect 1135 -754 1235 -554
rect 1293 -754 1393 -554
rect 1451 -754 1551 -554
rect 1609 -754 1709 -554
rect 1767 -754 1867 -554
rect 1925 -754 2025 -554
rect 2083 -754 2183 -554
rect -2183 -1190 -2083 -990
rect -2025 -1190 -1925 -990
rect -1867 -1190 -1767 -990
rect -1709 -1190 -1609 -990
rect -1551 -1190 -1451 -990
rect -1393 -1190 -1293 -990
rect -1235 -1190 -1135 -990
rect -1077 -1190 -977 -990
rect -919 -1190 -819 -990
rect -761 -1190 -661 -990
rect -603 -1190 -503 -990
rect -445 -1190 -345 -990
rect -287 -1190 -187 -990
rect -129 -1190 -29 -990
rect 29 -1190 129 -990
rect 187 -1190 287 -990
rect 345 -1190 445 -990
rect 503 -1190 603 -990
rect 661 -1190 761 -990
rect 819 -1190 919 -990
rect 977 -1190 1077 -990
rect 1135 -1190 1235 -990
rect 1293 -1190 1393 -990
rect 1451 -1190 1551 -990
rect 1609 -1190 1709 -990
rect 1767 -1190 1867 -990
rect 1925 -1190 2025 -990
rect 2083 -1190 2183 -990
rect -2183 -1626 -2083 -1426
rect -2025 -1626 -1925 -1426
rect -1867 -1626 -1767 -1426
rect -1709 -1626 -1609 -1426
rect -1551 -1626 -1451 -1426
rect -1393 -1626 -1293 -1426
rect -1235 -1626 -1135 -1426
rect -1077 -1626 -977 -1426
rect -919 -1626 -819 -1426
rect -761 -1626 -661 -1426
rect -603 -1626 -503 -1426
rect -445 -1626 -345 -1426
rect -287 -1626 -187 -1426
rect -129 -1626 -29 -1426
rect 29 -1626 129 -1426
rect 187 -1626 287 -1426
rect 345 -1626 445 -1426
rect 503 -1626 603 -1426
rect 661 -1626 761 -1426
rect 819 -1626 919 -1426
rect 977 -1626 1077 -1426
rect 1135 -1626 1235 -1426
rect 1293 -1626 1393 -1426
rect 1451 -1626 1551 -1426
rect 1609 -1626 1709 -1426
rect 1767 -1626 1867 -1426
rect 1925 -1626 2025 -1426
rect 2083 -1626 2183 -1426
rect -2183 -2062 -2083 -1862
rect -2025 -2062 -1925 -1862
rect -1867 -2062 -1767 -1862
rect -1709 -2062 -1609 -1862
rect -1551 -2062 -1451 -1862
rect -1393 -2062 -1293 -1862
rect -1235 -2062 -1135 -1862
rect -1077 -2062 -977 -1862
rect -919 -2062 -819 -1862
rect -761 -2062 -661 -1862
rect -603 -2062 -503 -1862
rect -445 -2062 -345 -1862
rect -287 -2062 -187 -1862
rect -129 -2062 -29 -1862
rect 29 -2062 129 -1862
rect 187 -2062 287 -1862
rect 345 -2062 445 -1862
rect 503 -2062 603 -1862
rect 661 -2062 761 -1862
rect 819 -2062 919 -1862
rect 977 -2062 1077 -1862
rect 1135 -2062 1235 -1862
rect 1293 -2062 1393 -1862
rect 1451 -2062 1551 -1862
rect 1609 -2062 1709 -1862
rect 1767 -2062 1867 -1862
rect 1925 -2062 2025 -1862
rect 2083 -2062 2183 -1862
<< mvpdiff >>
rect -2241 2050 -2183 2062
rect -2241 1874 -2229 2050
rect -2195 1874 -2183 2050
rect -2241 1862 -2183 1874
rect -2083 2050 -2025 2062
rect -2083 1874 -2071 2050
rect -2037 1874 -2025 2050
rect -2083 1862 -2025 1874
rect -1925 2050 -1867 2062
rect -1925 1874 -1913 2050
rect -1879 1874 -1867 2050
rect -1925 1862 -1867 1874
rect -1767 2050 -1709 2062
rect -1767 1874 -1755 2050
rect -1721 1874 -1709 2050
rect -1767 1862 -1709 1874
rect -1609 2050 -1551 2062
rect -1609 1874 -1597 2050
rect -1563 1874 -1551 2050
rect -1609 1862 -1551 1874
rect -1451 2050 -1393 2062
rect -1451 1874 -1439 2050
rect -1405 1874 -1393 2050
rect -1451 1862 -1393 1874
rect -1293 2050 -1235 2062
rect -1293 1874 -1281 2050
rect -1247 1874 -1235 2050
rect -1293 1862 -1235 1874
rect -1135 2050 -1077 2062
rect -1135 1874 -1123 2050
rect -1089 1874 -1077 2050
rect -1135 1862 -1077 1874
rect -977 2050 -919 2062
rect -977 1874 -965 2050
rect -931 1874 -919 2050
rect -977 1862 -919 1874
rect -819 2050 -761 2062
rect -819 1874 -807 2050
rect -773 1874 -761 2050
rect -819 1862 -761 1874
rect -661 2050 -603 2062
rect -661 1874 -649 2050
rect -615 1874 -603 2050
rect -661 1862 -603 1874
rect -503 2050 -445 2062
rect -503 1874 -491 2050
rect -457 1874 -445 2050
rect -503 1862 -445 1874
rect -345 2050 -287 2062
rect -345 1874 -333 2050
rect -299 1874 -287 2050
rect -345 1862 -287 1874
rect -187 2050 -129 2062
rect -187 1874 -175 2050
rect -141 1874 -129 2050
rect -187 1862 -129 1874
rect -29 2050 29 2062
rect -29 1874 -17 2050
rect 17 1874 29 2050
rect -29 1862 29 1874
rect 129 2050 187 2062
rect 129 1874 141 2050
rect 175 1874 187 2050
rect 129 1862 187 1874
rect 287 2050 345 2062
rect 287 1874 299 2050
rect 333 1874 345 2050
rect 287 1862 345 1874
rect 445 2050 503 2062
rect 445 1874 457 2050
rect 491 1874 503 2050
rect 445 1862 503 1874
rect 603 2050 661 2062
rect 603 1874 615 2050
rect 649 1874 661 2050
rect 603 1862 661 1874
rect 761 2050 819 2062
rect 761 1874 773 2050
rect 807 1874 819 2050
rect 761 1862 819 1874
rect 919 2050 977 2062
rect 919 1874 931 2050
rect 965 1874 977 2050
rect 919 1862 977 1874
rect 1077 2050 1135 2062
rect 1077 1874 1089 2050
rect 1123 1874 1135 2050
rect 1077 1862 1135 1874
rect 1235 2050 1293 2062
rect 1235 1874 1247 2050
rect 1281 1874 1293 2050
rect 1235 1862 1293 1874
rect 1393 2050 1451 2062
rect 1393 1874 1405 2050
rect 1439 1874 1451 2050
rect 1393 1862 1451 1874
rect 1551 2050 1609 2062
rect 1551 1874 1563 2050
rect 1597 1874 1609 2050
rect 1551 1862 1609 1874
rect 1709 2050 1767 2062
rect 1709 1874 1721 2050
rect 1755 1874 1767 2050
rect 1709 1862 1767 1874
rect 1867 2050 1925 2062
rect 1867 1874 1879 2050
rect 1913 1874 1925 2050
rect 1867 1862 1925 1874
rect 2025 2050 2083 2062
rect 2025 1874 2037 2050
rect 2071 1874 2083 2050
rect 2025 1862 2083 1874
rect 2183 2050 2241 2062
rect 2183 1874 2195 2050
rect 2229 1874 2241 2050
rect 2183 1862 2241 1874
rect -2241 1614 -2183 1626
rect -2241 1438 -2229 1614
rect -2195 1438 -2183 1614
rect -2241 1426 -2183 1438
rect -2083 1614 -2025 1626
rect -2083 1438 -2071 1614
rect -2037 1438 -2025 1614
rect -2083 1426 -2025 1438
rect -1925 1614 -1867 1626
rect -1925 1438 -1913 1614
rect -1879 1438 -1867 1614
rect -1925 1426 -1867 1438
rect -1767 1614 -1709 1626
rect -1767 1438 -1755 1614
rect -1721 1438 -1709 1614
rect -1767 1426 -1709 1438
rect -1609 1614 -1551 1626
rect -1609 1438 -1597 1614
rect -1563 1438 -1551 1614
rect -1609 1426 -1551 1438
rect -1451 1614 -1393 1626
rect -1451 1438 -1439 1614
rect -1405 1438 -1393 1614
rect -1451 1426 -1393 1438
rect -1293 1614 -1235 1626
rect -1293 1438 -1281 1614
rect -1247 1438 -1235 1614
rect -1293 1426 -1235 1438
rect -1135 1614 -1077 1626
rect -1135 1438 -1123 1614
rect -1089 1438 -1077 1614
rect -1135 1426 -1077 1438
rect -977 1614 -919 1626
rect -977 1438 -965 1614
rect -931 1438 -919 1614
rect -977 1426 -919 1438
rect -819 1614 -761 1626
rect -819 1438 -807 1614
rect -773 1438 -761 1614
rect -819 1426 -761 1438
rect -661 1614 -603 1626
rect -661 1438 -649 1614
rect -615 1438 -603 1614
rect -661 1426 -603 1438
rect -503 1614 -445 1626
rect -503 1438 -491 1614
rect -457 1438 -445 1614
rect -503 1426 -445 1438
rect -345 1614 -287 1626
rect -345 1438 -333 1614
rect -299 1438 -287 1614
rect -345 1426 -287 1438
rect -187 1614 -129 1626
rect -187 1438 -175 1614
rect -141 1438 -129 1614
rect -187 1426 -129 1438
rect -29 1614 29 1626
rect -29 1438 -17 1614
rect 17 1438 29 1614
rect -29 1426 29 1438
rect 129 1614 187 1626
rect 129 1438 141 1614
rect 175 1438 187 1614
rect 129 1426 187 1438
rect 287 1614 345 1626
rect 287 1438 299 1614
rect 333 1438 345 1614
rect 287 1426 345 1438
rect 445 1614 503 1626
rect 445 1438 457 1614
rect 491 1438 503 1614
rect 445 1426 503 1438
rect 603 1614 661 1626
rect 603 1438 615 1614
rect 649 1438 661 1614
rect 603 1426 661 1438
rect 761 1614 819 1626
rect 761 1438 773 1614
rect 807 1438 819 1614
rect 761 1426 819 1438
rect 919 1614 977 1626
rect 919 1438 931 1614
rect 965 1438 977 1614
rect 919 1426 977 1438
rect 1077 1614 1135 1626
rect 1077 1438 1089 1614
rect 1123 1438 1135 1614
rect 1077 1426 1135 1438
rect 1235 1614 1293 1626
rect 1235 1438 1247 1614
rect 1281 1438 1293 1614
rect 1235 1426 1293 1438
rect 1393 1614 1451 1626
rect 1393 1438 1405 1614
rect 1439 1438 1451 1614
rect 1393 1426 1451 1438
rect 1551 1614 1609 1626
rect 1551 1438 1563 1614
rect 1597 1438 1609 1614
rect 1551 1426 1609 1438
rect 1709 1614 1767 1626
rect 1709 1438 1721 1614
rect 1755 1438 1767 1614
rect 1709 1426 1767 1438
rect 1867 1614 1925 1626
rect 1867 1438 1879 1614
rect 1913 1438 1925 1614
rect 1867 1426 1925 1438
rect 2025 1614 2083 1626
rect 2025 1438 2037 1614
rect 2071 1438 2083 1614
rect 2025 1426 2083 1438
rect 2183 1614 2241 1626
rect 2183 1438 2195 1614
rect 2229 1438 2241 1614
rect 2183 1426 2241 1438
rect -2241 1178 -2183 1190
rect -2241 1002 -2229 1178
rect -2195 1002 -2183 1178
rect -2241 990 -2183 1002
rect -2083 1178 -2025 1190
rect -2083 1002 -2071 1178
rect -2037 1002 -2025 1178
rect -2083 990 -2025 1002
rect -1925 1178 -1867 1190
rect -1925 1002 -1913 1178
rect -1879 1002 -1867 1178
rect -1925 990 -1867 1002
rect -1767 1178 -1709 1190
rect -1767 1002 -1755 1178
rect -1721 1002 -1709 1178
rect -1767 990 -1709 1002
rect -1609 1178 -1551 1190
rect -1609 1002 -1597 1178
rect -1563 1002 -1551 1178
rect -1609 990 -1551 1002
rect -1451 1178 -1393 1190
rect -1451 1002 -1439 1178
rect -1405 1002 -1393 1178
rect -1451 990 -1393 1002
rect -1293 1178 -1235 1190
rect -1293 1002 -1281 1178
rect -1247 1002 -1235 1178
rect -1293 990 -1235 1002
rect -1135 1178 -1077 1190
rect -1135 1002 -1123 1178
rect -1089 1002 -1077 1178
rect -1135 990 -1077 1002
rect -977 1178 -919 1190
rect -977 1002 -965 1178
rect -931 1002 -919 1178
rect -977 990 -919 1002
rect -819 1178 -761 1190
rect -819 1002 -807 1178
rect -773 1002 -761 1178
rect -819 990 -761 1002
rect -661 1178 -603 1190
rect -661 1002 -649 1178
rect -615 1002 -603 1178
rect -661 990 -603 1002
rect -503 1178 -445 1190
rect -503 1002 -491 1178
rect -457 1002 -445 1178
rect -503 990 -445 1002
rect -345 1178 -287 1190
rect -345 1002 -333 1178
rect -299 1002 -287 1178
rect -345 990 -287 1002
rect -187 1178 -129 1190
rect -187 1002 -175 1178
rect -141 1002 -129 1178
rect -187 990 -129 1002
rect -29 1178 29 1190
rect -29 1002 -17 1178
rect 17 1002 29 1178
rect -29 990 29 1002
rect 129 1178 187 1190
rect 129 1002 141 1178
rect 175 1002 187 1178
rect 129 990 187 1002
rect 287 1178 345 1190
rect 287 1002 299 1178
rect 333 1002 345 1178
rect 287 990 345 1002
rect 445 1178 503 1190
rect 445 1002 457 1178
rect 491 1002 503 1178
rect 445 990 503 1002
rect 603 1178 661 1190
rect 603 1002 615 1178
rect 649 1002 661 1178
rect 603 990 661 1002
rect 761 1178 819 1190
rect 761 1002 773 1178
rect 807 1002 819 1178
rect 761 990 819 1002
rect 919 1178 977 1190
rect 919 1002 931 1178
rect 965 1002 977 1178
rect 919 990 977 1002
rect 1077 1178 1135 1190
rect 1077 1002 1089 1178
rect 1123 1002 1135 1178
rect 1077 990 1135 1002
rect 1235 1178 1293 1190
rect 1235 1002 1247 1178
rect 1281 1002 1293 1178
rect 1235 990 1293 1002
rect 1393 1178 1451 1190
rect 1393 1002 1405 1178
rect 1439 1002 1451 1178
rect 1393 990 1451 1002
rect 1551 1178 1609 1190
rect 1551 1002 1563 1178
rect 1597 1002 1609 1178
rect 1551 990 1609 1002
rect 1709 1178 1767 1190
rect 1709 1002 1721 1178
rect 1755 1002 1767 1178
rect 1709 990 1767 1002
rect 1867 1178 1925 1190
rect 1867 1002 1879 1178
rect 1913 1002 1925 1178
rect 1867 990 1925 1002
rect 2025 1178 2083 1190
rect 2025 1002 2037 1178
rect 2071 1002 2083 1178
rect 2025 990 2083 1002
rect 2183 1178 2241 1190
rect 2183 1002 2195 1178
rect 2229 1002 2241 1178
rect 2183 990 2241 1002
rect -2241 742 -2183 754
rect -2241 566 -2229 742
rect -2195 566 -2183 742
rect -2241 554 -2183 566
rect -2083 742 -2025 754
rect -2083 566 -2071 742
rect -2037 566 -2025 742
rect -2083 554 -2025 566
rect -1925 742 -1867 754
rect -1925 566 -1913 742
rect -1879 566 -1867 742
rect -1925 554 -1867 566
rect -1767 742 -1709 754
rect -1767 566 -1755 742
rect -1721 566 -1709 742
rect -1767 554 -1709 566
rect -1609 742 -1551 754
rect -1609 566 -1597 742
rect -1563 566 -1551 742
rect -1609 554 -1551 566
rect -1451 742 -1393 754
rect -1451 566 -1439 742
rect -1405 566 -1393 742
rect -1451 554 -1393 566
rect -1293 742 -1235 754
rect -1293 566 -1281 742
rect -1247 566 -1235 742
rect -1293 554 -1235 566
rect -1135 742 -1077 754
rect -1135 566 -1123 742
rect -1089 566 -1077 742
rect -1135 554 -1077 566
rect -977 742 -919 754
rect -977 566 -965 742
rect -931 566 -919 742
rect -977 554 -919 566
rect -819 742 -761 754
rect -819 566 -807 742
rect -773 566 -761 742
rect -819 554 -761 566
rect -661 742 -603 754
rect -661 566 -649 742
rect -615 566 -603 742
rect -661 554 -603 566
rect -503 742 -445 754
rect -503 566 -491 742
rect -457 566 -445 742
rect -503 554 -445 566
rect -345 742 -287 754
rect -345 566 -333 742
rect -299 566 -287 742
rect -345 554 -287 566
rect -187 742 -129 754
rect -187 566 -175 742
rect -141 566 -129 742
rect -187 554 -129 566
rect -29 742 29 754
rect -29 566 -17 742
rect 17 566 29 742
rect -29 554 29 566
rect 129 742 187 754
rect 129 566 141 742
rect 175 566 187 742
rect 129 554 187 566
rect 287 742 345 754
rect 287 566 299 742
rect 333 566 345 742
rect 287 554 345 566
rect 445 742 503 754
rect 445 566 457 742
rect 491 566 503 742
rect 445 554 503 566
rect 603 742 661 754
rect 603 566 615 742
rect 649 566 661 742
rect 603 554 661 566
rect 761 742 819 754
rect 761 566 773 742
rect 807 566 819 742
rect 761 554 819 566
rect 919 742 977 754
rect 919 566 931 742
rect 965 566 977 742
rect 919 554 977 566
rect 1077 742 1135 754
rect 1077 566 1089 742
rect 1123 566 1135 742
rect 1077 554 1135 566
rect 1235 742 1293 754
rect 1235 566 1247 742
rect 1281 566 1293 742
rect 1235 554 1293 566
rect 1393 742 1451 754
rect 1393 566 1405 742
rect 1439 566 1451 742
rect 1393 554 1451 566
rect 1551 742 1609 754
rect 1551 566 1563 742
rect 1597 566 1609 742
rect 1551 554 1609 566
rect 1709 742 1767 754
rect 1709 566 1721 742
rect 1755 566 1767 742
rect 1709 554 1767 566
rect 1867 742 1925 754
rect 1867 566 1879 742
rect 1913 566 1925 742
rect 1867 554 1925 566
rect 2025 742 2083 754
rect 2025 566 2037 742
rect 2071 566 2083 742
rect 2025 554 2083 566
rect 2183 742 2241 754
rect 2183 566 2195 742
rect 2229 566 2241 742
rect 2183 554 2241 566
rect -2241 306 -2183 318
rect -2241 130 -2229 306
rect -2195 130 -2183 306
rect -2241 118 -2183 130
rect -2083 306 -2025 318
rect -2083 130 -2071 306
rect -2037 130 -2025 306
rect -2083 118 -2025 130
rect -1925 306 -1867 318
rect -1925 130 -1913 306
rect -1879 130 -1867 306
rect -1925 118 -1867 130
rect -1767 306 -1709 318
rect -1767 130 -1755 306
rect -1721 130 -1709 306
rect -1767 118 -1709 130
rect -1609 306 -1551 318
rect -1609 130 -1597 306
rect -1563 130 -1551 306
rect -1609 118 -1551 130
rect -1451 306 -1393 318
rect -1451 130 -1439 306
rect -1405 130 -1393 306
rect -1451 118 -1393 130
rect -1293 306 -1235 318
rect -1293 130 -1281 306
rect -1247 130 -1235 306
rect -1293 118 -1235 130
rect -1135 306 -1077 318
rect -1135 130 -1123 306
rect -1089 130 -1077 306
rect -1135 118 -1077 130
rect -977 306 -919 318
rect -977 130 -965 306
rect -931 130 -919 306
rect -977 118 -919 130
rect -819 306 -761 318
rect -819 130 -807 306
rect -773 130 -761 306
rect -819 118 -761 130
rect -661 306 -603 318
rect -661 130 -649 306
rect -615 130 -603 306
rect -661 118 -603 130
rect -503 306 -445 318
rect -503 130 -491 306
rect -457 130 -445 306
rect -503 118 -445 130
rect -345 306 -287 318
rect -345 130 -333 306
rect -299 130 -287 306
rect -345 118 -287 130
rect -187 306 -129 318
rect -187 130 -175 306
rect -141 130 -129 306
rect -187 118 -129 130
rect -29 306 29 318
rect -29 130 -17 306
rect 17 130 29 306
rect -29 118 29 130
rect 129 306 187 318
rect 129 130 141 306
rect 175 130 187 306
rect 129 118 187 130
rect 287 306 345 318
rect 287 130 299 306
rect 333 130 345 306
rect 287 118 345 130
rect 445 306 503 318
rect 445 130 457 306
rect 491 130 503 306
rect 445 118 503 130
rect 603 306 661 318
rect 603 130 615 306
rect 649 130 661 306
rect 603 118 661 130
rect 761 306 819 318
rect 761 130 773 306
rect 807 130 819 306
rect 761 118 819 130
rect 919 306 977 318
rect 919 130 931 306
rect 965 130 977 306
rect 919 118 977 130
rect 1077 306 1135 318
rect 1077 130 1089 306
rect 1123 130 1135 306
rect 1077 118 1135 130
rect 1235 306 1293 318
rect 1235 130 1247 306
rect 1281 130 1293 306
rect 1235 118 1293 130
rect 1393 306 1451 318
rect 1393 130 1405 306
rect 1439 130 1451 306
rect 1393 118 1451 130
rect 1551 306 1609 318
rect 1551 130 1563 306
rect 1597 130 1609 306
rect 1551 118 1609 130
rect 1709 306 1767 318
rect 1709 130 1721 306
rect 1755 130 1767 306
rect 1709 118 1767 130
rect 1867 306 1925 318
rect 1867 130 1879 306
rect 1913 130 1925 306
rect 1867 118 1925 130
rect 2025 306 2083 318
rect 2025 130 2037 306
rect 2071 130 2083 306
rect 2025 118 2083 130
rect 2183 306 2241 318
rect 2183 130 2195 306
rect 2229 130 2241 306
rect 2183 118 2241 130
rect -2241 -130 -2183 -118
rect -2241 -306 -2229 -130
rect -2195 -306 -2183 -130
rect -2241 -318 -2183 -306
rect -2083 -130 -2025 -118
rect -2083 -306 -2071 -130
rect -2037 -306 -2025 -130
rect -2083 -318 -2025 -306
rect -1925 -130 -1867 -118
rect -1925 -306 -1913 -130
rect -1879 -306 -1867 -130
rect -1925 -318 -1867 -306
rect -1767 -130 -1709 -118
rect -1767 -306 -1755 -130
rect -1721 -306 -1709 -130
rect -1767 -318 -1709 -306
rect -1609 -130 -1551 -118
rect -1609 -306 -1597 -130
rect -1563 -306 -1551 -130
rect -1609 -318 -1551 -306
rect -1451 -130 -1393 -118
rect -1451 -306 -1439 -130
rect -1405 -306 -1393 -130
rect -1451 -318 -1393 -306
rect -1293 -130 -1235 -118
rect -1293 -306 -1281 -130
rect -1247 -306 -1235 -130
rect -1293 -318 -1235 -306
rect -1135 -130 -1077 -118
rect -1135 -306 -1123 -130
rect -1089 -306 -1077 -130
rect -1135 -318 -1077 -306
rect -977 -130 -919 -118
rect -977 -306 -965 -130
rect -931 -306 -919 -130
rect -977 -318 -919 -306
rect -819 -130 -761 -118
rect -819 -306 -807 -130
rect -773 -306 -761 -130
rect -819 -318 -761 -306
rect -661 -130 -603 -118
rect -661 -306 -649 -130
rect -615 -306 -603 -130
rect -661 -318 -603 -306
rect -503 -130 -445 -118
rect -503 -306 -491 -130
rect -457 -306 -445 -130
rect -503 -318 -445 -306
rect -345 -130 -287 -118
rect -345 -306 -333 -130
rect -299 -306 -287 -130
rect -345 -318 -287 -306
rect -187 -130 -129 -118
rect -187 -306 -175 -130
rect -141 -306 -129 -130
rect -187 -318 -129 -306
rect -29 -130 29 -118
rect -29 -306 -17 -130
rect 17 -306 29 -130
rect -29 -318 29 -306
rect 129 -130 187 -118
rect 129 -306 141 -130
rect 175 -306 187 -130
rect 129 -318 187 -306
rect 287 -130 345 -118
rect 287 -306 299 -130
rect 333 -306 345 -130
rect 287 -318 345 -306
rect 445 -130 503 -118
rect 445 -306 457 -130
rect 491 -306 503 -130
rect 445 -318 503 -306
rect 603 -130 661 -118
rect 603 -306 615 -130
rect 649 -306 661 -130
rect 603 -318 661 -306
rect 761 -130 819 -118
rect 761 -306 773 -130
rect 807 -306 819 -130
rect 761 -318 819 -306
rect 919 -130 977 -118
rect 919 -306 931 -130
rect 965 -306 977 -130
rect 919 -318 977 -306
rect 1077 -130 1135 -118
rect 1077 -306 1089 -130
rect 1123 -306 1135 -130
rect 1077 -318 1135 -306
rect 1235 -130 1293 -118
rect 1235 -306 1247 -130
rect 1281 -306 1293 -130
rect 1235 -318 1293 -306
rect 1393 -130 1451 -118
rect 1393 -306 1405 -130
rect 1439 -306 1451 -130
rect 1393 -318 1451 -306
rect 1551 -130 1609 -118
rect 1551 -306 1563 -130
rect 1597 -306 1609 -130
rect 1551 -318 1609 -306
rect 1709 -130 1767 -118
rect 1709 -306 1721 -130
rect 1755 -306 1767 -130
rect 1709 -318 1767 -306
rect 1867 -130 1925 -118
rect 1867 -306 1879 -130
rect 1913 -306 1925 -130
rect 1867 -318 1925 -306
rect 2025 -130 2083 -118
rect 2025 -306 2037 -130
rect 2071 -306 2083 -130
rect 2025 -318 2083 -306
rect 2183 -130 2241 -118
rect 2183 -306 2195 -130
rect 2229 -306 2241 -130
rect 2183 -318 2241 -306
rect -2241 -566 -2183 -554
rect -2241 -742 -2229 -566
rect -2195 -742 -2183 -566
rect -2241 -754 -2183 -742
rect -2083 -566 -2025 -554
rect -2083 -742 -2071 -566
rect -2037 -742 -2025 -566
rect -2083 -754 -2025 -742
rect -1925 -566 -1867 -554
rect -1925 -742 -1913 -566
rect -1879 -742 -1867 -566
rect -1925 -754 -1867 -742
rect -1767 -566 -1709 -554
rect -1767 -742 -1755 -566
rect -1721 -742 -1709 -566
rect -1767 -754 -1709 -742
rect -1609 -566 -1551 -554
rect -1609 -742 -1597 -566
rect -1563 -742 -1551 -566
rect -1609 -754 -1551 -742
rect -1451 -566 -1393 -554
rect -1451 -742 -1439 -566
rect -1405 -742 -1393 -566
rect -1451 -754 -1393 -742
rect -1293 -566 -1235 -554
rect -1293 -742 -1281 -566
rect -1247 -742 -1235 -566
rect -1293 -754 -1235 -742
rect -1135 -566 -1077 -554
rect -1135 -742 -1123 -566
rect -1089 -742 -1077 -566
rect -1135 -754 -1077 -742
rect -977 -566 -919 -554
rect -977 -742 -965 -566
rect -931 -742 -919 -566
rect -977 -754 -919 -742
rect -819 -566 -761 -554
rect -819 -742 -807 -566
rect -773 -742 -761 -566
rect -819 -754 -761 -742
rect -661 -566 -603 -554
rect -661 -742 -649 -566
rect -615 -742 -603 -566
rect -661 -754 -603 -742
rect -503 -566 -445 -554
rect -503 -742 -491 -566
rect -457 -742 -445 -566
rect -503 -754 -445 -742
rect -345 -566 -287 -554
rect -345 -742 -333 -566
rect -299 -742 -287 -566
rect -345 -754 -287 -742
rect -187 -566 -129 -554
rect -187 -742 -175 -566
rect -141 -742 -129 -566
rect -187 -754 -129 -742
rect -29 -566 29 -554
rect -29 -742 -17 -566
rect 17 -742 29 -566
rect -29 -754 29 -742
rect 129 -566 187 -554
rect 129 -742 141 -566
rect 175 -742 187 -566
rect 129 -754 187 -742
rect 287 -566 345 -554
rect 287 -742 299 -566
rect 333 -742 345 -566
rect 287 -754 345 -742
rect 445 -566 503 -554
rect 445 -742 457 -566
rect 491 -742 503 -566
rect 445 -754 503 -742
rect 603 -566 661 -554
rect 603 -742 615 -566
rect 649 -742 661 -566
rect 603 -754 661 -742
rect 761 -566 819 -554
rect 761 -742 773 -566
rect 807 -742 819 -566
rect 761 -754 819 -742
rect 919 -566 977 -554
rect 919 -742 931 -566
rect 965 -742 977 -566
rect 919 -754 977 -742
rect 1077 -566 1135 -554
rect 1077 -742 1089 -566
rect 1123 -742 1135 -566
rect 1077 -754 1135 -742
rect 1235 -566 1293 -554
rect 1235 -742 1247 -566
rect 1281 -742 1293 -566
rect 1235 -754 1293 -742
rect 1393 -566 1451 -554
rect 1393 -742 1405 -566
rect 1439 -742 1451 -566
rect 1393 -754 1451 -742
rect 1551 -566 1609 -554
rect 1551 -742 1563 -566
rect 1597 -742 1609 -566
rect 1551 -754 1609 -742
rect 1709 -566 1767 -554
rect 1709 -742 1721 -566
rect 1755 -742 1767 -566
rect 1709 -754 1767 -742
rect 1867 -566 1925 -554
rect 1867 -742 1879 -566
rect 1913 -742 1925 -566
rect 1867 -754 1925 -742
rect 2025 -566 2083 -554
rect 2025 -742 2037 -566
rect 2071 -742 2083 -566
rect 2025 -754 2083 -742
rect 2183 -566 2241 -554
rect 2183 -742 2195 -566
rect 2229 -742 2241 -566
rect 2183 -754 2241 -742
rect -2241 -1002 -2183 -990
rect -2241 -1178 -2229 -1002
rect -2195 -1178 -2183 -1002
rect -2241 -1190 -2183 -1178
rect -2083 -1002 -2025 -990
rect -2083 -1178 -2071 -1002
rect -2037 -1178 -2025 -1002
rect -2083 -1190 -2025 -1178
rect -1925 -1002 -1867 -990
rect -1925 -1178 -1913 -1002
rect -1879 -1178 -1867 -1002
rect -1925 -1190 -1867 -1178
rect -1767 -1002 -1709 -990
rect -1767 -1178 -1755 -1002
rect -1721 -1178 -1709 -1002
rect -1767 -1190 -1709 -1178
rect -1609 -1002 -1551 -990
rect -1609 -1178 -1597 -1002
rect -1563 -1178 -1551 -1002
rect -1609 -1190 -1551 -1178
rect -1451 -1002 -1393 -990
rect -1451 -1178 -1439 -1002
rect -1405 -1178 -1393 -1002
rect -1451 -1190 -1393 -1178
rect -1293 -1002 -1235 -990
rect -1293 -1178 -1281 -1002
rect -1247 -1178 -1235 -1002
rect -1293 -1190 -1235 -1178
rect -1135 -1002 -1077 -990
rect -1135 -1178 -1123 -1002
rect -1089 -1178 -1077 -1002
rect -1135 -1190 -1077 -1178
rect -977 -1002 -919 -990
rect -977 -1178 -965 -1002
rect -931 -1178 -919 -1002
rect -977 -1190 -919 -1178
rect -819 -1002 -761 -990
rect -819 -1178 -807 -1002
rect -773 -1178 -761 -1002
rect -819 -1190 -761 -1178
rect -661 -1002 -603 -990
rect -661 -1178 -649 -1002
rect -615 -1178 -603 -1002
rect -661 -1190 -603 -1178
rect -503 -1002 -445 -990
rect -503 -1178 -491 -1002
rect -457 -1178 -445 -1002
rect -503 -1190 -445 -1178
rect -345 -1002 -287 -990
rect -345 -1178 -333 -1002
rect -299 -1178 -287 -1002
rect -345 -1190 -287 -1178
rect -187 -1002 -129 -990
rect -187 -1178 -175 -1002
rect -141 -1178 -129 -1002
rect -187 -1190 -129 -1178
rect -29 -1002 29 -990
rect -29 -1178 -17 -1002
rect 17 -1178 29 -1002
rect -29 -1190 29 -1178
rect 129 -1002 187 -990
rect 129 -1178 141 -1002
rect 175 -1178 187 -1002
rect 129 -1190 187 -1178
rect 287 -1002 345 -990
rect 287 -1178 299 -1002
rect 333 -1178 345 -1002
rect 287 -1190 345 -1178
rect 445 -1002 503 -990
rect 445 -1178 457 -1002
rect 491 -1178 503 -1002
rect 445 -1190 503 -1178
rect 603 -1002 661 -990
rect 603 -1178 615 -1002
rect 649 -1178 661 -1002
rect 603 -1190 661 -1178
rect 761 -1002 819 -990
rect 761 -1178 773 -1002
rect 807 -1178 819 -1002
rect 761 -1190 819 -1178
rect 919 -1002 977 -990
rect 919 -1178 931 -1002
rect 965 -1178 977 -1002
rect 919 -1190 977 -1178
rect 1077 -1002 1135 -990
rect 1077 -1178 1089 -1002
rect 1123 -1178 1135 -1002
rect 1077 -1190 1135 -1178
rect 1235 -1002 1293 -990
rect 1235 -1178 1247 -1002
rect 1281 -1178 1293 -1002
rect 1235 -1190 1293 -1178
rect 1393 -1002 1451 -990
rect 1393 -1178 1405 -1002
rect 1439 -1178 1451 -1002
rect 1393 -1190 1451 -1178
rect 1551 -1002 1609 -990
rect 1551 -1178 1563 -1002
rect 1597 -1178 1609 -1002
rect 1551 -1190 1609 -1178
rect 1709 -1002 1767 -990
rect 1709 -1178 1721 -1002
rect 1755 -1178 1767 -1002
rect 1709 -1190 1767 -1178
rect 1867 -1002 1925 -990
rect 1867 -1178 1879 -1002
rect 1913 -1178 1925 -1002
rect 1867 -1190 1925 -1178
rect 2025 -1002 2083 -990
rect 2025 -1178 2037 -1002
rect 2071 -1178 2083 -1002
rect 2025 -1190 2083 -1178
rect 2183 -1002 2241 -990
rect 2183 -1178 2195 -1002
rect 2229 -1178 2241 -1002
rect 2183 -1190 2241 -1178
rect -2241 -1438 -2183 -1426
rect -2241 -1614 -2229 -1438
rect -2195 -1614 -2183 -1438
rect -2241 -1626 -2183 -1614
rect -2083 -1438 -2025 -1426
rect -2083 -1614 -2071 -1438
rect -2037 -1614 -2025 -1438
rect -2083 -1626 -2025 -1614
rect -1925 -1438 -1867 -1426
rect -1925 -1614 -1913 -1438
rect -1879 -1614 -1867 -1438
rect -1925 -1626 -1867 -1614
rect -1767 -1438 -1709 -1426
rect -1767 -1614 -1755 -1438
rect -1721 -1614 -1709 -1438
rect -1767 -1626 -1709 -1614
rect -1609 -1438 -1551 -1426
rect -1609 -1614 -1597 -1438
rect -1563 -1614 -1551 -1438
rect -1609 -1626 -1551 -1614
rect -1451 -1438 -1393 -1426
rect -1451 -1614 -1439 -1438
rect -1405 -1614 -1393 -1438
rect -1451 -1626 -1393 -1614
rect -1293 -1438 -1235 -1426
rect -1293 -1614 -1281 -1438
rect -1247 -1614 -1235 -1438
rect -1293 -1626 -1235 -1614
rect -1135 -1438 -1077 -1426
rect -1135 -1614 -1123 -1438
rect -1089 -1614 -1077 -1438
rect -1135 -1626 -1077 -1614
rect -977 -1438 -919 -1426
rect -977 -1614 -965 -1438
rect -931 -1614 -919 -1438
rect -977 -1626 -919 -1614
rect -819 -1438 -761 -1426
rect -819 -1614 -807 -1438
rect -773 -1614 -761 -1438
rect -819 -1626 -761 -1614
rect -661 -1438 -603 -1426
rect -661 -1614 -649 -1438
rect -615 -1614 -603 -1438
rect -661 -1626 -603 -1614
rect -503 -1438 -445 -1426
rect -503 -1614 -491 -1438
rect -457 -1614 -445 -1438
rect -503 -1626 -445 -1614
rect -345 -1438 -287 -1426
rect -345 -1614 -333 -1438
rect -299 -1614 -287 -1438
rect -345 -1626 -287 -1614
rect -187 -1438 -129 -1426
rect -187 -1614 -175 -1438
rect -141 -1614 -129 -1438
rect -187 -1626 -129 -1614
rect -29 -1438 29 -1426
rect -29 -1614 -17 -1438
rect 17 -1614 29 -1438
rect -29 -1626 29 -1614
rect 129 -1438 187 -1426
rect 129 -1614 141 -1438
rect 175 -1614 187 -1438
rect 129 -1626 187 -1614
rect 287 -1438 345 -1426
rect 287 -1614 299 -1438
rect 333 -1614 345 -1438
rect 287 -1626 345 -1614
rect 445 -1438 503 -1426
rect 445 -1614 457 -1438
rect 491 -1614 503 -1438
rect 445 -1626 503 -1614
rect 603 -1438 661 -1426
rect 603 -1614 615 -1438
rect 649 -1614 661 -1438
rect 603 -1626 661 -1614
rect 761 -1438 819 -1426
rect 761 -1614 773 -1438
rect 807 -1614 819 -1438
rect 761 -1626 819 -1614
rect 919 -1438 977 -1426
rect 919 -1614 931 -1438
rect 965 -1614 977 -1438
rect 919 -1626 977 -1614
rect 1077 -1438 1135 -1426
rect 1077 -1614 1089 -1438
rect 1123 -1614 1135 -1438
rect 1077 -1626 1135 -1614
rect 1235 -1438 1293 -1426
rect 1235 -1614 1247 -1438
rect 1281 -1614 1293 -1438
rect 1235 -1626 1293 -1614
rect 1393 -1438 1451 -1426
rect 1393 -1614 1405 -1438
rect 1439 -1614 1451 -1438
rect 1393 -1626 1451 -1614
rect 1551 -1438 1609 -1426
rect 1551 -1614 1563 -1438
rect 1597 -1614 1609 -1438
rect 1551 -1626 1609 -1614
rect 1709 -1438 1767 -1426
rect 1709 -1614 1721 -1438
rect 1755 -1614 1767 -1438
rect 1709 -1626 1767 -1614
rect 1867 -1438 1925 -1426
rect 1867 -1614 1879 -1438
rect 1913 -1614 1925 -1438
rect 1867 -1626 1925 -1614
rect 2025 -1438 2083 -1426
rect 2025 -1614 2037 -1438
rect 2071 -1614 2083 -1438
rect 2025 -1626 2083 -1614
rect 2183 -1438 2241 -1426
rect 2183 -1614 2195 -1438
rect 2229 -1614 2241 -1438
rect 2183 -1626 2241 -1614
rect -2241 -1874 -2183 -1862
rect -2241 -2050 -2229 -1874
rect -2195 -2050 -2183 -1874
rect -2241 -2062 -2183 -2050
rect -2083 -1874 -2025 -1862
rect -2083 -2050 -2071 -1874
rect -2037 -2050 -2025 -1874
rect -2083 -2062 -2025 -2050
rect -1925 -1874 -1867 -1862
rect -1925 -2050 -1913 -1874
rect -1879 -2050 -1867 -1874
rect -1925 -2062 -1867 -2050
rect -1767 -1874 -1709 -1862
rect -1767 -2050 -1755 -1874
rect -1721 -2050 -1709 -1874
rect -1767 -2062 -1709 -2050
rect -1609 -1874 -1551 -1862
rect -1609 -2050 -1597 -1874
rect -1563 -2050 -1551 -1874
rect -1609 -2062 -1551 -2050
rect -1451 -1874 -1393 -1862
rect -1451 -2050 -1439 -1874
rect -1405 -2050 -1393 -1874
rect -1451 -2062 -1393 -2050
rect -1293 -1874 -1235 -1862
rect -1293 -2050 -1281 -1874
rect -1247 -2050 -1235 -1874
rect -1293 -2062 -1235 -2050
rect -1135 -1874 -1077 -1862
rect -1135 -2050 -1123 -1874
rect -1089 -2050 -1077 -1874
rect -1135 -2062 -1077 -2050
rect -977 -1874 -919 -1862
rect -977 -2050 -965 -1874
rect -931 -2050 -919 -1874
rect -977 -2062 -919 -2050
rect -819 -1874 -761 -1862
rect -819 -2050 -807 -1874
rect -773 -2050 -761 -1874
rect -819 -2062 -761 -2050
rect -661 -1874 -603 -1862
rect -661 -2050 -649 -1874
rect -615 -2050 -603 -1874
rect -661 -2062 -603 -2050
rect -503 -1874 -445 -1862
rect -503 -2050 -491 -1874
rect -457 -2050 -445 -1874
rect -503 -2062 -445 -2050
rect -345 -1874 -287 -1862
rect -345 -2050 -333 -1874
rect -299 -2050 -287 -1874
rect -345 -2062 -287 -2050
rect -187 -1874 -129 -1862
rect -187 -2050 -175 -1874
rect -141 -2050 -129 -1874
rect -187 -2062 -129 -2050
rect -29 -1874 29 -1862
rect -29 -2050 -17 -1874
rect 17 -2050 29 -1874
rect -29 -2062 29 -2050
rect 129 -1874 187 -1862
rect 129 -2050 141 -1874
rect 175 -2050 187 -1874
rect 129 -2062 187 -2050
rect 287 -1874 345 -1862
rect 287 -2050 299 -1874
rect 333 -2050 345 -1874
rect 287 -2062 345 -2050
rect 445 -1874 503 -1862
rect 445 -2050 457 -1874
rect 491 -2050 503 -1874
rect 445 -2062 503 -2050
rect 603 -1874 661 -1862
rect 603 -2050 615 -1874
rect 649 -2050 661 -1874
rect 603 -2062 661 -2050
rect 761 -1874 819 -1862
rect 761 -2050 773 -1874
rect 807 -2050 819 -1874
rect 761 -2062 819 -2050
rect 919 -1874 977 -1862
rect 919 -2050 931 -1874
rect 965 -2050 977 -1874
rect 919 -2062 977 -2050
rect 1077 -1874 1135 -1862
rect 1077 -2050 1089 -1874
rect 1123 -2050 1135 -1874
rect 1077 -2062 1135 -2050
rect 1235 -1874 1293 -1862
rect 1235 -2050 1247 -1874
rect 1281 -2050 1293 -1874
rect 1235 -2062 1293 -2050
rect 1393 -1874 1451 -1862
rect 1393 -2050 1405 -1874
rect 1439 -2050 1451 -1874
rect 1393 -2062 1451 -2050
rect 1551 -1874 1609 -1862
rect 1551 -2050 1563 -1874
rect 1597 -2050 1609 -1874
rect 1551 -2062 1609 -2050
rect 1709 -1874 1767 -1862
rect 1709 -2050 1721 -1874
rect 1755 -2050 1767 -1874
rect 1709 -2062 1767 -2050
rect 1867 -1874 1925 -1862
rect 1867 -2050 1879 -1874
rect 1913 -2050 1925 -1874
rect 1867 -2062 1925 -2050
rect 2025 -1874 2083 -1862
rect 2025 -2050 2037 -1874
rect 2071 -2050 2083 -1874
rect 2025 -2062 2083 -2050
rect 2183 -1874 2241 -1862
rect 2183 -2050 2195 -1874
rect 2229 -2050 2241 -1874
rect 2183 -2062 2241 -2050
<< mvpdiffc >>
rect -2229 1874 -2195 2050
rect -2071 1874 -2037 2050
rect -1913 1874 -1879 2050
rect -1755 1874 -1721 2050
rect -1597 1874 -1563 2050
rect -1439 1874 -1405 2050
rect -1281 1874 -1247 2050
rect -1123 1874 -1089 2050
rect -965 1874 -931 2050
rect -807 1874 -773 2050
rect -649 1874 -615 2050
rect -491 1874 -457 2050
rect -333 1874 -299 2050
rect -175 1874 -141 2050
rect -17 1874 17 2050
rect 141 1874 175 2050
rect 299 1874 333 2050
rect 457 1874 491 2050
rect 615 1874 649 2050
rect 773 1874 807 2050
rect 931 1874 965 2050
rect 1089 1874 1123 2050
rect 1247 1874 1281 2050
rect 1405 1874 1439 2050
rect 1563 1874 1597 2050
rect 1721 1874 1755 2050
rect 1879 1874 1913 2050
rect 2037 1874 2071 2050
rect 2195 1874 2229 2050
rect -2229 1438 -2195 1614
rect -2071 1438 -2037 1614
rect -1913 1438 -1879 1614
rect -1755 1438 -1721 1614
rect -1597 1438 -1563 1614
rect -1439 1438 -1405 1614
rect -1281 1438 -1247 1614
rect -1123 1438 -1089 1614
rect -965 1438 -931 1614
rect -807 1438 -773 1614
rect -649 1438 -615 1614
rect -491 1438 -457 1614
rect -333 1438 -299 1614
rect -175 1438 -141 1614
rect -17 1438 17 1614
rect 141 1438 175 1614
rect 299 1438 333 1614
rect 457 1438 491 1614
rect 615 1438 649 1614
rect 773 1438 807 1614
rect 931 1438 965 1614
rect 1089 1438 1123 1614
rect 1247 1438 1281 1614
rect 1405 1438 1439 1614
rect 1563 1438 1597 1614
rect 1721 1438 1755 1614
rect 1879 1438 1913 1614
rect 2037 1438 2071 1614
rect 2195 1438 2229 1614
rect -2229 1002 -2195 1178
rect -2071 1002 -2037 1178
rect -1913 1002 -1879 1178
rect -1755 1002 -1721 1178
rect -1597 1002 -1563 1178
rect -1439 1002 -1405 1178
rect -1281 1002 -1247 1178
rect -1123 1002 -1089 1178
rect -965 1002 -931 1178
rect -807 1002 -773 1178
rect -649 1002 -615 1178
rect -491 1002 -457 1178
rect -333 1002 -299 1178
rect -175 1002 -141 1178
rect -17 1002 17 1178
rect 141 1002 175 1178
rect 299 1002 333 1178
rect 457 1002 491 1178
rect 615 1002 649 1178
rect 773 1002 807 1178
rect 931 1002 965 1178
rect 1089 1002 1123 1178
rect 1247 1002 1281 1178
rect 1405 1002 1439 1178
rect 1563 1002 1597 1178
rect 1721 1002 1755 1178
rect 1879 1002 1913 1178
rect 2037 1002 2071 1178
rect 2195 1002 2229 1178
rect -2229 566 -2195 742
rect -2071 566 -2037 742
rect -1913 566 -1879 742
rect -1755 566 -1721 742
rect -1597 566 -1563 742
rect -1439 566 -1405 742
rect -1281 566 -1247 742
rect -1123 566 -1089 742
rect -965 566 -931 742
rect -807 566 -773 742
rect -649 566 -615 742
rect -491 566 -457 742
rect -333 566 -299 742
rect -175 566 -141 742
rect -17 566 17 742
rect 141 566 175 742
rect 299 566 333 742
rect 457 566 491 742
rect 615 566 649 742
rect 773 566 807 742
rect 931 566 965 742
rect 1089 566 1123 742
rect 1247 566 1281 742
rect 1405 566 1439 742
rect 1563 566 1597 742
rect 1721 566 1755 742
rect 1879 566 1913 742
rect 2037 566 2071 742
rect 2195 566 2229 742
rect -2229 130 -2195 306
rect -2071 130 -2037 306
rect -1913 130 -1879 306
rect -1755 130 -1721 306
rect -1597 130 -1563 306
rect -1439 130 -1405 306
rect -1281 130 -1247 306
rect -1123 130 -1089 306
rect -965 130 -931 306
rect -807 130 -773 306
rect -649 130 -615 306
rect -491 130 -457 306
rect -333 130 -299 306
rect -175 130 -141 306
rect -17 130 17 306
rect 141 130 175 306
rect 299 130 333 306
rect 457 130 491 306
rect 615 130 649 306
rect 773 130 807 306
rect 931 130 965 306
rect 1089 130 1123 306
rect 1247 130 1281 306
rect 1405 130 1439 306
rect 1563 130 1597 306
rect 1721 130 1755 306
rect 1879 130 1913 306
rect 2037 130 2071 306
rect 2195 130 2229 306
rect -2229 -306 -2195 -130
rect -2071 -306 -2037 -130
rect -1913 -306 -1879 -130
rect -1755 -306 -1721 -130
rect -1597 -306 -1563 -130
rect -1439 -306 -1405 -130
rect -1281 -306 -1247 -130
rect -1123 -306 -1089 -130
rect -965 -306 -931 -130
rect -807 -306 -773 -130
rect -649 -306 -615 -130
rect -491 -306 -457 -130
rect -333 -306 -299 -130
rect -175 -306 -141 -130
rect -17 -306 17 -130
rect 141 -306 175 -130
rect 299 -306 333 -130
rect 457 -306 491 -130
rect 615 -306 649 -130
rect 773 -306 807 -130
rect 931 -306 965 -130
rect 1089 -306 1123 -130
rect 1247 -306 1281 -130
rect 1405 -306 1439 -130
rect 1563 -306 1597 -130
rect 1721 -306 1755 -130
rect 1879 -306 1913 -130
rect 2037 -306 2071 -130
rect 2195 -306 2229 -130
rect -2229 -742 -2195 -566
rect -2071 -742 -2037 -566
rect -1913 -742 -1879 -566
rect -1755 -742 -1721 -566
rect -1597 -742 -1563 -566
rect -1439 -742 -1405 -566
rect -1281 -742 -1247 -566
rect -1123 -742 -1089 -566
rect -965 -742 -931 -566
rect -807 -742 -773 -566
rect -649 -742 -615 -566
rect -491 -742 -457 -566
rect -333 -742 -299 -566
rect -175 -742 -141 -566
rect -17 -742 17 -566
rect 141 -742 175 -566
rect 299 -742 333 -566
rect 457 -742 491 -566
rect 615 -742 649 -566
rect 773 -742 807 -566
rect 931 -742 965 -566
rect 1089 -742 1123 -566
rect 1247 -742 1281 -566
rect 1405 -742 1439 -566
rect 1563 -742 1597 -566
rect 1721 -742 1755 -566
rect 1879 -742 1913 -566
rect 2037 -742 2071 -566
rect 2195 -742 2229 -566
rect -2229 -1178 -2195 -1002
rect -2071 -1178 -2037 -1002
rect -1913 -1178 -1879 -1002
rect -1755 -1178 -1721 -1002
rect -1597 -1178 -1563 -1002
rect -1439 -1178 -1405 -1002
rect -1281 -1178 -1247 -1002
rect -1123 -1178 -1089 -1002
rect -965 -1178 -931 -1002
rect -807 -1178 -773 -1002
rect -649 -1178 -615 -1002
rect -491 -1178 -457 -1002
rect -333 -1178 -299 -1002
rect -175 -1178 -141 -1002
rect -17 -1178 17 -1002
rect 141 -1178 175 -1002
rect 299 -1178 333 -1002
rect 457 -1178 491 -1002
rect 615 -1178 649 -1002
rect 773 -1178 807 -1002
rect 931 -1178 965 -1002
rect 1089 -1178 1123 -1002
rect 1247 -1178 1281 -1002
rect 1405 -1178 1439 -1002
rect 1563 -1178 1597 -1002
rect 1721 -1178 1755 -1002
rect 1879 -1178 1913 -1002
rect 2037 -1178 2071 -1002
rect 2195 -1178 2229 -1002
rect -2229 -1614 -2195 -1438
rect -2071 -1614 -2037 -1438
rect -1913 -1614 -1879 -1438
rect -1755 -1614 -1721 -1438
rect -1597 -1614 -1563 -1438
rect -1439 -1614 -1405 -1438
rect -1281 -1614 -1247 -1438
rect -1123 -1614 -1089 -1438
rect -965 -1614 -931 -1438
rect -807 -1614 -773 -1438
rect -649 -1614 -615 -1438
rect -491 -1614 -457 -1438
rect -333 -1614 -299 -1438
rect -175 -1614 -141 -1438
rect -17 -1614 17 -1438
rect 141 -1614 175 -1438
rect 299 -1614 333 -1438
rect 457 -1614 491 -1438
rect 615 -1614 649 -1438
rect 773 -1614 807 -1438
rect 931 -1614 965 -1438
rect 1089 -1614 1123 -1438
rect 1247 -1614 1281 -1438
rect 1405 -1614 1439 -1438
rect 1563 -1614 1597 -1438
rect 1721 -1614 1755 -1438
rect 1879 -1614 1913 -1438
rect 2037 -1614 2071 -1438
rect 2195 -1614 2229 -1438
rect -2229 -2050 -2195 -1874
rect -2071 -2050 -2037 -1874
rect -1913 -2050 -1879 -1874
rect -1755 -2050 -1721 -1874
rect -1597 -2050 -1563 -1874
rect -1439 -2050 -1405 -1874
rect -1281 -2050 -1247 -1874
rect -1123 -2050 -1089 -1874
rect -965 -2050 -931 -1874
rect -807 -2050 -773 -1874
rect -649 -2050 -615 -1874
rect -491 -2050 -457 -1874
rect -333 -2050 -299 -1874
rect -175 -2050 -141 -1874
rect -17 -2050 17 -1874
rect 141 -2050 175 -1874
rect 299 -2050 333 -1874
rect 457 -2050 491 -1874
rect 615 -2050 649 -1874
rect 773 -2050 807 -1874
rect 931 -2050 965 -1874
rect 1089 -2050 1123 -1874
rect 1247 -2050 1281 -1874
rect 1405 -2050 1439 -1874
rect 1563 -2050 1597 -1874
rect 1721 -2050 1755 -1874
rect 1879 -2050 1913 -1874
rect 2037 -2050 2071 -1874
rect 2195 -2050 2229 -1874
<< mvnsubdiff >>
rect -2375 2281 2375 2293
rect -2375 2247 -2267 2281
rect 2267 2247 2375 2281
rect -2375 2235 2375 2247
rect -2375 2185 -2317 2235
rect -2375 -2185 -2363 2185
rect -2329 -2185 -2317 2185
rect 2317 2185 2375 2235
rect -2375 -2235 -2317 -2185
rect 2317 -2185 2329 2185
rect 2363 -2185 2375 2185
rect 2317 -2235 2375 -2185
rect -2375 -2247 2375 -2235
rect -2375 -2281 -2267 -2247
rect 2267 -2281 2375 -2247
rect -2375 -2293 2375 -2281
<< mvnsubdiffcont >>
rect -2267 2247 2267 2281
rect -2363 -2185 -2329 2185
rect 2329 -2185 2363 2185
rect -2267 -2281 2267 -2247
<< poly >>
rect -2183 2143 -2083 2159
rect -2183 2109 -2167 2143
rect -2099 2109 -2083 2143
rect -2183 2062 -2083 2109
rect -2025 2143 -1925 2159
rect -2025 2109 -2009 2143
rect -1941 2109 -1925 2143
rect -2025 2062 -1925 2109
rect -1867 2143 -1767 2159
rect -1867 2109 -1851 2143
rect -1783 2109 -1767 2143
rect -1867 2062 -1767 2109
rect -1709 2143 -1609 2159
rect -1709 2109 -1693 2143
rect -1625 2109 -1609 2143
rect -1709 2062 -1609 2109
rect -1551 2143 -1451 2159
rect -1551 2109 -1535 2143
rect -1467 2109 -1451 2143
rect -1551 2062 -1451 2109
rect -1393 2143 -1293 2159
rect -1393 2109 -1377 2143
rect -1309 2109 -1293 2143
rect -1393 2062 -1293 2109
rect -1235 2143 -1135 2159
rect -1235 2109 -1219 2143
rect -1151 2109 -1135 2143
rect -1235 2062 -1135 2109
rect -1077 2143 -977 2159
rect -1077 2109 -1061 2143
rect -993 2109 -977 2143
rect -1077 2062 -977 2109
rect -919 2143 -819 2159
rect -919 2109 -903 2143
rect -835 2109 -819 2143
rect -919 2062 -819 2109
rect -761 2143 -661 2159
rect -761 2109 -745 2143
rect -677 2109 -661 2143
rect -761 2062 -661 2109
rect -603 2143 -503 2159
rect -603 2109 -587 2143
rect -519 2109 -503 2143
rect -603 2062 -503 2109
rect -445 2143 -345 2159
rect -445 2109 -429 2143
rect -361 2109 -345 2143
rect -445 2062 -345 2109
rect -287 2143 -187 2159
rect -287 2109 -271 2143
rect -203 2109 -187 2143
rect -287 2062 -187 2109
rect -129 2143 -29 2159
rect -129 2109 -113 2143
rect -45 2109 -29 2143
rect -129 2062 -29 2109
rect 29 2143 129 2159
rect 29 2109 45 2143
rect 113 2109 129 2143
rect 29 2062 129 2109
rect 187 2143 287 2159
rect 187 2109 203 2143
rect 271 2109 287 2143
rect 187 2062 287 2109
rect 345 2143 445 2159
rect 345 2109 361 2143
rect 429 2109 445 2143
rect 345 2062 445 2109
rect 503 2143 603 2159
rect 503 2109 519 2143
rect 587 2109 603 2143
rect 503 2062 603 2109
rect 661 2143 761 2159
rect 661 2109 677 2143
rect 745 2109 761 2143
rect 661 2062 761 2109
rect 819 2143 919 2159
rect 819 2109 835 2143
rect 903 2109 919 2143
rect 819 2062 919 2109
rect 977 2143 1077 2159
rect 977 2109 993 2143
rect 1061 2109 1077 2143
rect 977 2062 1077 2109
rect 1135 2143 1235 2159
rect 1135 2109 1151 2143
rect 1219 2109 1235 2143
rect 1135 2062 1235 2109
rect 1293 2143 1393 2159
rect 1293 2109 1309 2143
rect 1377 2109 1393 2143
rect 1293 2062 1393 2109
rect 1451 2143 1551 2159
rect 1451 2109 1467 2143
rect 1535 2109 1551 2143
rect 1451 2062 1551 2109
rect 1609 2143 1709 2159
rect 1609 2109 1625 2143
rect 1693 2109 1709 2143
rect 1609 2062 1709 2109
rect 1767 2143 1867 2159
rect 1767 2109 1783 2143
rect 1851 2109 1867 2143
rect 1767 2062 1867 2109
rect 1925 2143 2025 2159
rect 1925 2109 1941 2143
rect 2009 2109 2025 2143
rect 1925 2062 2025 2109
rect 2083 2143 2183 2159
rect 2083 2109 2099 2143
rect 2167 2109 2183 2143
rect 2083 2062 2183 2109
rect -2183 1815 -2083 1862
rect -2183 1781 -2167 1815
rect -2099 1781 -2083 1815
rect -2183 1765 -2083 1781
rect -2025 1815 -1925 1862
rect -2025 1781 -2009 1815
rect -1941 1781 -1925 1815
rect -2025 1765 -1925 1781
rect -1867 1815 -1767 1862
rect -1867 1781 -1851 1815
rect -1783 1781 -1767 1815
rect -1867 1765 -1767 1781
rect -1709 1815 -1609 1862
rect -1709 1781 -1693 1815
rect -1625 1781 -1609 1815
rect -1709 1765 -1609 1781
rect -1551 1815 -1451 1862
rect -1551 1781 -1535 1815
rect -1467 1781 -1451 1815
rect -1551 1765 -1451 1781
rect -1393 1815 -1293 1862
rect -1393 1781 -1377 1815
rect -1309 1781 -1293 1815
rect -1393 1765 -1293 1781
rect -1235 1815 -1135 1862
rect -1235 1781 -1219 1815
rect -1151 1781 -1135 1815
rect -1235 1765 -1135 1781
rect -1077 1815 -977 1862
rect -1077 1781 -1061 1815
rect -993 1781 -977 1815
rect -1077 1765 -977 1781
rect -919 1815 -819 1862
rect -919 1781 -903 1815
rect -835 1781 -819 1815
rect -919 1765 -819 1781
rect -761 1815 -661 1862
rect -761 1781 -745 1815
rect -677 1781 -661 1815
rect -761 1765 -661 1781
rect -603 1815 -503 1862
rect -603 1781 -587 1815
rect -519 1781 -503 1815
rect -603 1765 -503 1781
rect -445 1815 -345 1862
rect -445 1781 -429 1815
rect -361 1781 -345 1815
rect -445 1765 -345 1781
rect -287 1815 -187 1862
rect -287 1781 -271 1815
rect -203 1781 -187 1815
rect -287 1765 -187 1781
rect -129 1815 -29 1862
rect -129 1781 -113 1815
rect -45 1781 -29 1815
rect -129 1765 -29 1781
rect 29 1815 129 1862
rect 29 1781 45 1815
rect 113 1781 129 1815
rect 29 1765 129 1781
rect 187 1815 287 1862
rect 187 1781 203 1815
rect 271 1781 287 1815
rect 187 1765 287 1781
rect 345 1815 445 1862
rect 345 1781 361 1815
rect 429 1781 445 1815
rect 345 1765 445 1781
rect 503 1815 603 1862
rect 503 1781 519 1815
rect 587 1781 603 1815
rect 503 1765 603 1781
rect 661 1815 761 1862
rect 661 1781 677 1815
rect 745 1781 761 1815
rect 661 1765 761 1781
rect 819 1815 919 1862
rect 819 1781 835 1815
rect 903 1781 919 1815
rect 819 1765 919 1781
rect 977 1815 1077 1862
rect 977 1781 993 1815
rect 1061 1781 1077 1815
rect 977 1765 1077 1781
rect 1135 1815 1235 1862
rect 1135 1781 1151 1815
rect 1219 1781 1235 1815
rect 1135 1765 1235 1781
rect 1293 1815 1393 1862
rect 1293 1781 1309 1815
rect 1377 1781 1393 1815
rect 1293 1765 1393 1781
rect 1451 1815 1551 1862
rect 1451 1781 1467 1815
rect 1535 1781 1551 1815
rect 1451 1765 1551 1781
rect 1609 1815 1709 1862
rect 1609 1781 1625 1815
rect 1693 1781 1709 1815
rect 1609 1765 1709 1781
rect 1767 1815 1867 1862
rect 1767 1781 1783 1815
rect 1851 1781 1867 1815
rect 1767 1765 1867 1781
rect 1925 1815 2025 1862
rect 1925 1781 1941 1815
rect 2009 1781 2025 1815
rect 1925 1765 2025 1781
rect 2083 1815 2183 1862
rect 2083 1781 2099 1815
rect 2167 1781 2183 1815
rect 2083 1765 2183 1781
rect -2183 1707 -2083 1723
rect -2183 1673 -2167 1707
rect -2099 1673 -2083 1707
rect -2183 1626 -2083 1673
rect -2025 1707 -1925 1723
rect -2025 1673 -2009 1707
rect -1941 1673 -1925 1707
rect -2025 1626 -1925 1673
rect -1867 1707 -1767 1723
rect -1867 1673 -1851 1707
rect -1783 1673 -1767 1707
rect -1867 1626 -1767 1673
rect -1709 1707 -1609 1723
rect -1709 1673 -1693 1707
rect -1625 1673 -1609 1707
rect -1709 1626 -1609 1673
rect -1551 1707 -1451 1723
rect -1551 1673 -1535 1707
rect -1467 1673 -1451 1707
rect -1551 1626 -1451 1673
rect -1393 1707 -1293 1723
rect -1393 1673 -1377 1707
rect -1309 1673 -1293 1707
rect -1393 1626 -1293 1673
rect -1235 1707 -1135 1723
rect -1235 1673 -1219 1707
rect -1151 1673 -1135 1707
rect -1235 1626 -1135 1673
rect -1077 1707 -977 1723
rect -1077 1673 -1061 1707
rect -993 1673 -977 1707
rect -1077 1626 -977 1673
rect -919 1707 -819 1723
rect -919 1673 -903 1707
rect -835 1673 -819 1707
rect -919 1626 -819 1673
rect -761 1707 -661 1723
rect -761 1673 -745 1707
rect -677 1673 -661 1707
rect -761 1626 -661 1673
rect -603 1707 -503 1723
rect -603 1673 -587 1707
rect -519 1673 -503 1707
rect -603 1626 -503 1673
rect -445 1707 -345 1723
rect -445 1673 -429 1707
rect -361 1673 -345 1707
rect -445 1626 -345 1673
rect -287 1707 -187 1723
rect -287 1673 -271 1707
rect -203 1673 -187 1707
rect -287 1626 -187 1673
rect -129 1707 -29 1723
rect -129 1673 -113 1707
rect -45 1673 -29 1707
rect -129 1626 -29 1673
rect 29 1707 129 1723
rect 29 1673 45 1707
rect 113 1673 129 1707
rect 29 1626 129 1673
rect 187 1707 287 1723
rect 187 1673 203 1707
rect 271 1673 287 1707
rect 187 1626 287 1673
rect 345 1707 445 1723
rect 345 1673 361 1707
rect 429 1673 445 1707
rect 345 1626 445 1673
rect 503 1707 603 1723
rect 503 1673 519 1707
rect 587 1673 603 1707
rect 503 1626 603 1673
rect 661 1707 761 1723
rect 661 1673 677 1707
rect 745 1673 761 1707
rect 661 1626 761 1673
rect 819 1707 919 1723
rect 819 1673 835 1707
rect 903 1673 919 1707
rect 819 1626 919 1673
rect 977 1707 1077 1723
rect 977 1673 993 1707
rect 1061 1673 1077 1707
rect 977 1626 1077 1673
rect 1135 1707 1235 1723
rect 1135 1673 1151 1707
rect 1219 1673 1235 1707
rect 1135 1626 1235 1673
rect 1293 1707 1393 1723
rect 1293 1673 1309 1707
rect 1377 1673 1393 1707
rect 1293 1626 1393 1673
rect 1451 1707 1551 1723
rect 1451 1673 1467 1707
rect 1535 1673 1551 1707
rect 1451 1626 1551 1673
rect 1609 1707 1709 1723
rect 1609 1673 1625 1707
rect 1693 1673 1709 1707
rect 1609 1626 1709 1673
rect 1767 1707 1867 1723
rect 1767 1673 1783 1707
rect 1851 1673 1867 1707
rect 1767 1626 1867 1673
rect 1925 1707 2025 1723
rect 1925 1673 1941 1707
rect 2009 1673 2025 1707
rect 1925 1626 2025 1673
rect 2083 1707 2183 1723
rect 2083 1673 2099 1707
rect 2167 1673 2183 1707
rect 2083 1626 2183 1673
rect -2183 1379 -2083 1426
rect -2183 1345 -2167 1379
rect -2099 1345 -2083 1379
rect -2183 1329 -2083 1345
rect -2025 1379 -1925 1426
rect -2025 1345 -2009 1379
rect -1941 1345 -1925 1379
rect -2025 1329 -1925 1345
rect -1867 1379 -1767 1426
rect -1867 1345 -1851 1379
rect -1783 1345 -1767 1379
rect -1867 1329 -1767 1345
rect -1709 1379 -1609 1426
rect -1709 1345 -1693 1379
rect -1625 1345 -1609 1379
rect -1709 1329 -1609 1345
rect -1551 1379 -1451 1426
rect -1551 1345 -1535 1379
rect -1467 1345 -1451 1379
rect -1551 1329 -1451 1345
rect -1393 1379 -1293 1426
rect -1393 1345 -1377 1379
rect -1309 1345 -1293 1379
rect -1393 1329 -1293 1345
rect -1235 1379 -1135 1426
rect -1235 1345 -1219 1379
rect -1151 1345 -1135 1379
rect -1235 1329 -1135 1345
rect -1077 1379 -977 1426
rect -1077 1345 -1061 1379
rect -993 1345 -977 1379
rect -1077 1329 -977 1345
rect -919 1379 -819 1426
rect -919 1345 -903 1379
rect -835 1345 -819 1379
rect -919 1329 -819 1345
rect -761 1379 -661 1426
rect -761 1345 -745 1379
rect -677 1345 -661 1379
rect -761 1329 -661 1345
rect -603 1379 -503 1426
rect -603 1345 -587 1379
rect -519 1345 -503 1379
rect -603 1329 -503 1345
rect -445 1379 -345 1426
rect -445 1345 -429 1379
rect -361 1345 -345 1379
rect -445 1329 -345 1345
rect -287 1379 -187 1426
rect -287 1345 -271 1379
rect -203 1345 -187 1379
rect -287 1329 -187 1345
rect -129 1379 -29 1426
rect -129 1345 -113 1379
rect -45 1345 -29 1379
rect -129 1329 -29 1345
rect 29 1379 129 1426
rect 29 1345 45 1379
rect 113 1345 129 1379
rect 29 1329 129 1345
rect 187 1379 287 1426
rect 187 1345 203 1379
rect 271 1345 287 1379
rect 187 1329 287 1345
rect 345 1379 445 1426
rect 345 1345 361 1379
rect 429 1345 445 1379
rect 345 1329 445 1345
rect 503 1379 603 1426
rect 503 1345 519 1379
rect 587 1345 603 1379
rect 503 1329 603 1345
rect 661 1379 761 1426
rect 661 1345 677 1379
rect 745 1345 761 1379
rect 661 1329 761 1345
rect 819 1379 919 1426
rect 819 1345 835 1379
rect 903 1345 919 1379
rect 819 1329 919 1345
rect 977 1379 1077 1426
rect 977 1345 993 1379
rect 1061 1345 1077 1379
rect 977 1329 1077 1345
rect 1135 1379 1235 1426
rect 1135 1345 1151 1379
rect 1219 1345 1235 1379
rect 1135 1329 1235 1345
rect 1293 1379 1393 1426
rect 1293 1345 1309 1379
rect 1377 1345 1393 1379
rect 1293 1329 1393 1345
rect 1451 1379 1551 1426
rect 1451 1345 1467 1379
rect 1535 1345 1551 1379
rect 1451 1329 1551 1345
rect 1609 1379 1709 1426
rect 1609 1345 1625 1379
rect 1693 1345 1709 1379
rect 1609 1329 1709 1345
rect 1767 1379 1867 1426
rect 1767 1345 1783 1379
rect 1851 1345 1867 1379
rect 1767 1329 1867 1345
rect 1925 1379 2025 1426
rect 1925 1345 1941 1379
rect 2009 1345 2025 1379
rect 1925 1329 2025 1345
rect 2083 1379 2183 1426
rect 2083 1345 2099 1379
rect 2167 1345 2183 1379
rect 2083 1329 2183 1345
rect -2183 1271 -2083 1287
rect -2183 1237 -2167 1271
rect -2099 1237 -2083 1271
rect -2183 1190 -2083 1237
rect -2025 1271 -1925 1287
rect -2025 1237 -2009 1271
rect -1941 1237 -1925 1271
rect -2025 1190 -1925 1237
rect -1867 1271 -1767 1287
rect -1867 1237 -1851 1271
rect -1783 1237 -1767 1271
rect -1867 1190 -1767 1237
rect -1709 1271 -1609 1287
rect -1709 1237 -1693 1271
rect -1625 1237 -1609 1271
rect -1709 1190 -1609 1237
rect -1551 1271 -1451 1287
rect -1551 1237 -1535 1271
rect -1467 1237 -1451 1271
rect -1551 1190 -1451 1237
rect -1393 1271 -1293 1287
rect -1393 1237 -1377 1271
rect -1309 1237 -1293 1271
rect -1393 1190 -1293 1237
rect -1235 1271 -1135 1287
rect -1235 1237 -1219 1271
rect -1151 1237 -1135 1271
rect -1235 1190 -1135 1237
rect -1077 1271 -977 1287
rect -1077 1237 -1061 1271
rect -993 1237 -977 1271
rect -1077 1190 -977 1237
rect -919 1271 -819 1287
rect -919 1237 -903 1271
rect -835 1237 -819 1271
rect -919 1190 -819 1237
rect -761 1271 -661 1287
rect -761 1237 -745 1271
rect -677 1237 -661 1271
rect -761 1190 -661 1237
rect -603 1271 -503 1287
rect -603 1237 -587 1271
rect -519 1237 -503 1271
rect -603 1190 -503 1237
rect -445 1271 -345 1287
rect -445 1237 -429 1271
rect -361 1237 -345 1271
rect -445 1190 -345 1237
rect -287 1271 -187 1287
rect -287 1237 -271 1271
rect -203 1237 -187 1271
rect -287 1190 -187 1237
rect -129 1271 -29 1287
rect -129 1237 -113 1271
rect -45 1237 -29 1271
rect -129 1190 -29 1237
rect 29 1271 129 1287
rect 29 1237 45 1271
rect 113 1237 129 1271
rect 29 1190 129 1237
rect 187 1271 287 1287
rect 187 1237 203 1271
rect 271 1237 287 1271
rect 187 1190 287 1237
rect 345 1271 445 1287
rect 345 1237 361 1271
rect 429 1237 445 1271
rect 345 1190 445 1237
rect 503 1271 603 1287
rect 503 1237 519 1271
rect 587 1237 603 1271
rect 503 1190 603 1237
rect 661 1271 761 1287
rect 661 1237 677 1271
rect 745 1237 761 1271
rect 661 1190 761 1237
rect 819 1271 919 1287
rect 819 1237 835 1271
rect 903 1237 919 1271
rect 819 1190 919 1237
rect 977 1271 1077 1287
rect 977 1237 993 1271
rect 1061 1237 1077 1271
rect 977 1190 1077 1237
rect 1135 1271 1235 1287
rect 1135 1237 1151 1271
rect 1219 1237 1235 1271
rect 1135 1190 1235 1237
rect 1293 1271 1393 1287
rect 1293 1237 1309 1271
rect 1377 1237 1393 1271
rect 1293 1190 1393 1237
rect 1451 1271 1551 1287
rect 1451 1237 1467 1271
rect 1535 1237 1551 1271
rect 1451 1190 1551 1237
rect 1609 1271 1709 1287
rect 1609 1237 1625 1271
rect 1693 1237 1709 1271
rect 1609 1190 1709 1237
rect 1767 1271 1867 1287
rect 1767 1237 1783 1271
rect 1851 1237 1867 1271
rect 1767 1190 1867 1237
rect 1925 1271 2025 1287
rect 1925 1237 1941 1271
rect 2009 1237 2025 1271
rect 1925 1190 2025 1237
rect 2083 1271 2183 1287
rect 2083 1237 2099 1271
rect 2167 1237 2183 1271
rect 2083 1190 2183 1237
rect -2183 943 -2083 990
rect -2183 909 -2167 943
rect -2099 909 -2083 943
rect -2183 893 -2083 909
rect -2025 943 -1925 990
rect -2025 909 -2009 943
rect -1941 909 -1925 943
rect -2025 893 -1925 909
rect -1867 943 -1767 990
rect -1867 909 -1851 943
rect -1783 909 -1767 943
rect -1867 893 -1767 909
rect -1709 943 -1609 990
rect -1709 909 -1693 943
rect -1625 909 -1609 943
rect -1709 893 -1609 909
rect -1551 943 -1451 990
rect -1551 909 -1535 943
rect -1467 909 -1451 943
rect -1551 893 -1451 909
rect -1393 943 -1293 990
rect -1393 909 -1377 943
rect -1309 909 -1293 943
rect -1393 893 -1293 909
rect -1235 943 -1135 990
rect -1235 909 -1219 943
rect -1151 909 -1135 943
rect -1235 893 -1135 909
rect -1077 943 -977 990
rect -1077 909 -1061 943
rect -993 909 -977 943
rect -1077 893 -977 909
rect -919 943 -819 990
rect -919 909 -903 943
rect -835 909 -819 943
rect -919 893 -819 909
rect -761 943 -661 990
rect -761 909 -745 943
rect -677 909 -661 943
rect -761 893 -661 909
rect -603 943 -503 990
rect -603 909 -587 943
rect -519 909 -503 943
rect -603 893 -503 909
rect -445 943 -345 990
rect -445 909 -429 943
rect -361 909 -345 943
rect -445 893 -345 909
rect -287 943 -187 990
rect -287 909 -271 943
rect -203 909 -187 943
rect -287 893 -187 909
rect -129 943 -29 990
rect -129 909 -113 943
rect -45 909 -29 943
rect -129 893 -29 909
rect 29 943 129 990
rect 29 909 45 943
rect 113 909 129 943
rect 29 893 129 909
rect 187 943 287 990
rect 187 909 203 943
rect 271 909 287 943
rect 187 893 287 909
rect 345 943 445 990
rect 345 909 361 943
rect 429 909 445 943
rect 345 893 445 909
rect 503 943 603 990
rect 503 909 519 943
rect 587 909 603 943
rect 503 893 603 909
rect 661 943 761 990
rect 661 909 677 943
rect 745 909 761 943
rect 661 893 761 909
rect 819 943 919 990
rect 819 909 835 943
rect 903 909 919 943
rect 819 893 919 909
rect 977 943 1077 990
rect 977 909 993 943
rect 1061 909 1077 943
rect 977 893 1077 909
rect 1135 943 1235 990
rect 1135 909 1151 943
rect 1219 909 1235 943
rect 1135 893 1235 909
rect 1293 943 1393 990
rect 1293 909 1309 943
rect 1377 909 1393 943
rect 1293 893 1393 909
rect 1451 943 1551 990
rect 1451 909 1467 943
rect 1535 909 1551 943
rect 1451 893 1551 909
rect 1609 943 1709 990
rect 1609 909 1625 943
rect 1693 909 1709 943
rect 1609 893 1709 909
rect 1767 943 1867 990
rect 1767 909 1783 943
rect 1851 909 1867 943
rect 1767 893 1867 909
rect 1925 943 2025 990
rect 1925 909 1941 943
rect 2009 909 2025 943
rect 1925 893 2025 909
rect 2083 943 2183 990
rect 2083 909 2099 943
rect 2167 909 2183 943
rect 2083 893 2183 909
rect -2183 835 -2083 851
rect -2183 801 -2167 835
rect -2099 801 -2083 835
rect -2183 754 -2083 801
rect -2025 835 -1925 851
rect -2025 801 -2009 835
rect -1941 801 -1925 835
rect -2025 754 -1925 801
rect -1867 835 -1767 851
rect -1867 801 -1851 835
rect -1783 801 -1767 835
rect -1867 754 -1767 801
rect -1709 835 -1609 851
rect -1709 801 -1693 835
rect -1625 801 -1609 835
rect -1709 754 -1609 801
rect -1551 835 -1451 851
rect -1551 801 -1535 835
rect -1467 801 -1451 835
rect -1551 754 -1451 801
rect -1393 835 -1293 851
rect -1393 801 -1377 835
rect -1309 801 -1293 835
rect -1393 754 -1293 801
rect -1235 835 -1135 851
rect -1235 801 -1219 835
rect -1151 801 -1135 835
rect -1235 754 -1135 801
rect -1077 835 -977 851
rect -1077 801 -1061 835
rect -993 801 -977 835
rect -1077 754 -977 801
rect -919 835 -819 851
rect -919 801 -903 835
rect -835 801 -819 835
rect -919 754 -819 801
rect -761 835 -661 851
rect -761 801 -745 835
rect -677 801 -661 835
rect -761 754 -661 801
rect -603 835 -503 851
rect -603 801 -587 835
rect -519 801 -503 835
rect -603 754 -503 801
rect -445 835 -345 851
rect -445 801 -429 835
rect -361 801 -345 835
rect -445 754 -345 801
rect -287 835 -187 851
rect -287 801 -271 835
rect -203 801 -187 835
rect -287 754 -187 801
rect -129 835 -29 851
rect -129 801 -113 835
rect -45 801 -29 835
rect -129 754 -29 801
rect 29 835 129 851
rect 29 801 45 835
rect 113 801 129 835
rect 29 754 129 801
rect 187 835 287 851
rect 187 801 203 835
rect 271 801 287 835
rect 187 754 287 801
rect 345 835 445 851
rect 345 801 361 835
rect 429 801 445 835
rect 345 754 445 801
rect 503 835 603 851
rect 503 801 519 835
rect 587 801 603 835
rect 503 754 603 801
rect 661 835 761 851
rect 661 801 677 835
rect 745 801 761 835
rect 661 754 761 801
rect 819 835 919 851
rect 819 801 835 835
rect 903 801 919 835
rect 819 754 919 801
rect 977 835 1077 851
rect 977 801 993 835
rect 1061 801 1077 835
rect 977 754 1077 801
rect 1135 835 1235 851
rect 1135 801 1151 835
rect 1219 801 1235 835
rect 1135 754 1235 801
rect 1293 835 1393 851
rect 1293 801 1309 835
rect 1377 801 1393 835
rect 1293 754 1393 801
rect 1451 835 1551 851
rect 1451 801 1467 835
rect 1535 801 1551 835
rect 1451 754 1551 801
rect 1609 835 1709 851
rect 1609 801 1625 835
rect 1693 801 1709 835
rect 1609 754 1709 801
rect 1767 835 1867 851
rect 1767 801 1783 835
rect 1851 801 1867 835
rect 1767 754 1867 801
rect 1925 835 2025 851
rect 1925 801 1941 835
rect 2009 801 2025 835
rect 1925 754 2025 801
rect 2083 835 2183 851
rect 2083 801 2099 835
rect 2167 801 2183 835
rect 2083 754 2183 801
rect -2183 507 -2083 554
rect -2183 473 -2167 507
rect -2099 473 -2083 507
rect -2183 457 -2083 473
rect -2025 507 -1925 554
rect -2025 473 -2009 507
rect -1941 473 -1925 507
rect -2025 457 -1925 473
rect -1867 507 -1767 554
rect -1867 473 -1851 507
rect -1783 473 -1767 507
rect -1867 457 -1767 473
rect -1709 507 -1609 554
rect -1709 473 -1693 507
rect -1625 473 -1609 507
rect -1709 457 -1609 473
rect -1551 507 -1451 554
rect -1551 473 -1535 507
rect -1467 473 -1451 507
rect -1551 457 -1451 473
rect -1393 507 -1293 554
rect -1393 473 -1377 507
rect -1309 473 -1293 507
rect -1393 457 -1293 473
rect -1235 507 -1135 554
rect -1235 473 -1219 507
rect -1151 473 -1135 507
rect -1235 457 -1135 473
rect -1077 507 -977 554
rect -1077 473 -1061 507
rect -993 473 -977 507
rect -1077 457 -977 473
rect -919 507 -819 554
rect -919 473 -903 507
rect -835 473 -819 507
rect -919 457 -819 473
rect -761 507 -661 554
rect -761 473 -745 507
rect -677 473 -661 507
rect -761 457 -661 473
rect -603 507 -503 554
rect -603 473 -587 507
rect -519 473 -503 507
rect -603 457 -503 473
rect -445 507 -345 554
rect -445 473 -429 507
rect -361 473 -345 507
rect -445 457 -345 473
rect -287 507 -187 554
rect -287 473 -271 507
rect -203 473 -187 507
rect -287 457 -187 473
rect -129 507 -29 554
rect -129 473 -113 507
rect -45 473 -29 507
rect -129 457 -29 473
rect 29 507 129 554
rect 29 473 45 507
rect 113 473 129 507
rect 29 457 129 473
rect 187 507 287 554
rect 187 473 203 507
rect 271 473 287 507
rect 187 457 287 473
rect 345 507 445 554
rect 345 473 361 507
rect 429 473 445 507
rect 345 457 445 473
rect 503 507 603 554
rect 503 473 519 507
rect 587 473 603 507
rect 503 457 603 473
rect 661 507 761 554
rect 661 473 677 507
rect 745 473 761 507
rect 661 457 761 473
rect 819 507 919 554
rect 819 473 835 507
rect 903 473 919 507
rect 819 457 919 473
rect 977 507 1077 554
rect 977 473 993 507
rect 1061 473 1077 507
rect 977 457 1077 473
rect 1135 507 1235 554
rect 1135 473 1151 507
rect 1219 473 1235 507
rect 1135 457 1235 473
rect 1293 507 1393 554
rect 1293 473 1309 507
rect 1377 473 1393 507
rect 1293 457 1393 473
rect 1451 507 1551 554
rect 1451 473 1467 507
rect 1535 473 1551 507
rect 1451 457 1551 473
rect 1609 507 1709 554
rect 1609 473 1625 507
rect 1693 473 1709 507
rect 1609 457 1709 473
rect 1767 507 1867 554
rect 1767 473 1783 507
rect 1851 473 1867 507
rect 1767 457 1867 473
rect 1925 507 2025 554
rect 1925 473 1941 507
rect 2009 473 2025 507
rect 1925 457 2025 473
rect 2083 507 2183 554
rect 2083 473 2099 507
rect 2167 473 2183 507
rect 2083 457 2183 473
rect -2183 399 -2083 415
rect -2183 365 -2167 399
rect -2099 365 -2083 399
rect -2183 318 -2083 365
rect -2025 399 -1925 415
rect -2025 365 -2009 399
rect -1941 365 -1925 399
rect -2025 318 -1925 365
rect -1867 399 -1767 415
rect -1867 365 -1851 399
rect -1783 365 -1767 399
rect -1867 318 -1767 365
rect -1709 399 -1609 415
rect -1709 365 -1693 399
rect -1625 365 -1609 399
rect -1709 318 -1609 365
rect -1551 399 -1451 415
rect -1551 365 -1535 399
rect -1467 365 -1451 399
rect -1551 318 -1451 365
rect -1393 399 -1293 415
rect -1393 365 -1377 399
rect -1309 365 -1293 399
rect -1393 318 -1293 365
rect -1235 399 -1135 415
rect -1235 365 -1219 399
rect -1151 365 -1135 399
rect -1235 318 -1135 365
rect -1077 399 -977 415
rect -1077 365 -1061 399
rect -993 365 -977 399
rect -1077 318 -977 365
rect -919 399 -819 415
rect -919 365 -903 399
rect -835 365 -819 399
rect -919 318 -819 365
rect -761 399 -661 415
rect -761 365 -745 399
rect -677 365 -661 399
rect -761 318 -661 365
rect -603 399 -503 415
rect -603 365 -587 399
rect -519 365 -503 399
rect -603 318 -503 365
rect -445 399 -345 415
rect -445 365 -429 399
rect -361 365 -345 399
rect -445 318 -345 365
rect -287 399 -187 415
rect -287 365 -271 399
rect -203 365 -187 399
rect -287 318 -187 365
rect -129 399 -29 415
rect -129 365 -113 399
rect -45 365 -29 399
rect -129 318 -29 365
rect 29 399 129 415
rect 29 365 45 399
rect 113 365 129 399
rect 29 318 129 365
rect 187 399 287 415
rect 187 365 203 399
rect 271 365 287 399
rect 187 318 287 365
rect 345 399 445 415
rect 345 365 361 399
rect 429 365 445 399
rect 345 318 445 365
rect 503 399 603 415
rect 503 365 519 399
rect 587 365 603 399
rect 503 318 603 365
rect 661 399 761 415
rect 661 365 677 399
rect 745 365 761 399
rect 661 318 761 365
rect 819 399 919 415
rect 819 365 835 399
rect 903 365 919 399
rect 819 318 919 365
rect 977 399 1077 415
rect 977 365 993 399
rect 1061 365 1077 399
rect 977 318 1077 365
rect 1135 399 1235 415
rect 1135 365 1151 399
rect 1219 365 1235 399
rect 1135 318 1235 365
rect 1293 399 1393 415
rect 1293 365 1309 399
rect 1377 365 1393 399
rect 1293 318 1393 365
rect 1451 399 1551 415
rect 1451 365 1467 399
rect 1535 365 1551 399
rect 1451 318 1551 365
rect 1609 399 1709 415
rect 1609 365 1625 399
rect 1693 365 1709 399
rect 1609 318 1709 365
rect 1767 399 1867 415
rect 1767 365 1783 399
rect 1851 365 1867 399
rect 1767 318 1867 365
rect 1925 399 2025 415
rect 1925 365 1941 399
rect 2009 365 2025 399
rect 1925 318 2025 365
rect 2083 399 2183 415
rect 2083 365 2099 399
rect 2167 365 2183 399
rect 2083 318 2183 365
rect -2183 71 -2083 118
rect -2183 37 -2167 71
rect -2099 37 -2083 71
rect -2183 21 -2083 37
rect -2025 71 -1925 118
rect -2025 37 -2009 71
rect -1941 37 -1925 71
rect -2025 21 -1925 37
rect -1867 71 -1767 118
rect -1867 37 -1851 71
rect -1783 37 -1767 71
rect -1867 21 -1767 37
rect -1709 71 -1609 118
rect -1709 37 -1693 71
rect -1625 37 -1609 71
rect -1709 21 -1609 37
rect -1551 71 -1451 118
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1551 21 -1451 37
rect -1393 71 -1293 118
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1393 21 -1293 37
rect -1235 71 -1135 118
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1235 21 -1135 37
rect -1077 71 -977 118
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -1077 21 -977 37
rect -919 71 -819 118
rect -919 37 -903 71
rect -835 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 118
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 118
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 118
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 118
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 118
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 118
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 118
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 118
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect 819 71 919 118
rect 819 37 835 71
rect 903 37 919 71
rect 819 21 919 37
rect 977 71 1077 118
rect 977 37 993 71
rect 1061 37 1077 71
rect 977 21 1077 37
rect 1135 71 1235 118
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1135 21 1235 37
rect 1293 71 1393 118
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1293 21 1393 37
rect 1451 71 1551 118
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1451 21 1551 37
rect 1609 71 1709 118
rect 1609 37 1625 71
rect 1693 37 1709 71
rect 1609 21 1709 37
rect 1767 71 1867 118
rect 1767 37 1783 71
rect 1851 37 1867 71
rect 1767 21 1867 37
rect 1925 71 2025 118
rect 1925 37 1941 71
rect 2009 37 2025 71
rect 1925 21 2025 37
rect 2083 71 2183 118
rect 2083 37 2099 71
rect 2167 37 2183 71
rect 2083 21 2183 37
rect -2183 -37 -2083 -21
rect -2183 -71 -2167 -37
rect -2099 -71 -2083 -37
rect -2183 -118 -2083 -71
rect -2025 -37 -1925 -21
rect -2025 -71 -2009 -37
rect -1941 -71 -1925 -37
rect -2025 -118 -1925 -71
rect -1867 -37 -1767 -21
rect -1867 -71 -1851 -37
rect -1783 -71 -1767 -37
rect -1867 -118 -1767 -71
rect -1709 -37 -1609 -21
rect -1709 -71 -1693 -37
rect -1625 -71 -1609 -37
rect -1709 -118 -1609 -71
rect -1551 -37 -1451 -21
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1551 -118 -1451 -71
rect -1393 -37 -1293 -21
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1393 -118 -1293 -71
rect -1235 -37 -1135 -21
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1235 -118 -1135 -71
rect -1077 -37 -977 -21
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -1077 -118 -977 -71
rect -919 -37 -819 -21
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -919 -118 -819 -71
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -118 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -118 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -118 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -118 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -118 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -118 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -118 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -118 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -118 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -118 761 -71
rect 819 -37 919 -21
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 819 -118 919 -71
rect 977 -37 1077 -21
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 977 -118 1077 -71
rect 1135 -37 1235 -21
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1135 -118 1235 -71
rect 1293 -37 1393 -21
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1293 -118 1393 -71
rect 1451 -37 1551 -21
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1451 -118 1551 -71
rect 1609 -37 1709 -21
rect 1609 -71 1625 -37
rect 1693 -71 1709 -37
rect 1609 -118 1709 -71
rect 1767 -37 1867 -21
rect 1767 -71 1783 -37
rect 1851 -71 1867 -37
rect 1767 -118 1867 -71
rect 1925 -37 2025 -21
rect 1925 -71 1941 -37
rect 2009 -71 2025 -37
rect 1925 -118 2025 -71
rect 2083 -37 2183 -21
rect 2083 -71 2099 -37
rect 2167 -71 2183 -37
rect 2083 -118 2183 -71
rect -2183 -365 -2083 -318
rect -2183 -399 -2167 -365
rect -2099 -399 -2083 -365
rect -2183 -415 -2083 -399
rect -2025 -365 -1925 -318
rect -2025 -399 -2009 -365
rect -1941 -399 -1925 -365
rect -2025 -415 -1925 -399
rect -1867 -365 -1767 -318
rect -1867 -399 -1851 -365
rect -1783 -399 -1767 -365
rect -1867 -415 -1767 -399
rect -1709 -365 -1609 -318
rect -1709 -399 -1693 -365
rect -1625 -399 -1609 -365
rect -1709 -415 -1609 -399
rect -1551 -365 -1451 -318
rect -1551 -399 -1535 -365
rect -1467 -399 -1451 -365
rect -1551 -415 -1451 -399
rect -1393 -365 -1293 -318
rect -1393 -399 -1377 -365
rect -1309 -399 -1293 -365
rect -1393 -415 -1293 -399
rect -1235 -365 -1135 -318
rect -1235 -399 -1219 -365
rect -1151 -399 -1135 -365
rect -1235 -415 -1135 -399
rect -1077 -365 -977 -318
rect -1077 -399 -1061 -365
rect -993 -399 -977 -365
rect -1077 -415 -977 -399
rect -919 -365 -819 -318
rect -919 -399 -903 -365
rect -835 -399 -819 -365
rect -919 -415 -819 -399
rect -761 -365 -661 -318
rect -761 -399 -745 -365
rect -677 -399 -661 -365
rect -761 -415 -661 -399
rect -603 -365 -503 -318
rect -603 -399 -587 -365
rect -519 -399 -503 -365
rect -603 -415 -503 -399
rect -445 -365 -345 -318
rect -445 -399 -429 -365
rect -361 -399 -345 -365
rect -445 -415 -345 -399
rect -287 -365 -187 -318
rect -287 -399 -271 -365
rect -203 -399 -187 -365
rect -287 -415 -187 -399
rect -129 -365 -29 -318
rect -129 -399 -113 -365
rect -45 -399 -29 -365
rect -129 -415 -29 -399
rect 29 -365 129 -318
rect 29 -399 45 -365
rect 113 -399 129 -365
rect 29 -415 129 -399
rect 187 -365 287 -318
rect 187 -399 203 -365
rect 271 -399 287 -365
rect 187 -415 287 -399
rect 345 -365 445 -318
rect 345 -399 361 -365
rect 429 -399 445 -365
rect 345 -415 445 -399
rect 503 -365 603 -318
rect 503 -399 519 -365
rect 587 -399 603 -365
rect 503 -415 603 -399
rect 661 -365 761 -318
rect 661 -399 677 -365
rect 745 -399 761 -365
rect 661 -415 761 -399
rect 819 -365 919 -318
rect 819 -399 835 -365
rect 903 -399 919 -365
rect 819 -415 919 -399
rect 977 -365 1077 -318
rect 977 -399 993 -365
rect 1061 -399 1077 -365
rect 977 -415 1077 -399
rect 1135 -365 1235 -318
rect 1135 -399 1151 -365
rect 1219 -399 1235 -365
rect 1135 -415 1235 -399
rect 1293 -365 1393 -318
rect 1293 -399 1309 -365
rect 1377 -399 1393 -365
rect 1293 -415 1393 -399
rect 1451 -365 1551 -318
rect 1451 -399 1467 -365
rect 1535 -399 1551 -365
rect 1451 -415 1551 -399
rect 1609 -365 1709 -318
rect 1609 -399 1625 -365
rect 1693 -399 1709 -365
rect 1609 -415 1709 -399
rect 1767 -365 1867 -318
rect 1767 -399 1783 -365
rect 1851 -399 1867 -365
rect 1767 -415 1867 -399
rect 1925 -365 2025 -318
rect 1925 -399 1941 -365
rect 2009 -399 2025 -365
rect 1925 -415 2025 -399
rect 2083 -365 2183 -318
rect 2083 -399 2099 -365
rect 2167 -399 2183 -365
rect 2083 -415 2183 -399
rect -2183 -473 -2083 -457
rect -2183 -507 -2167 -473
rect -2099 -507 -2083 -473
rect -2183 -554 -2083 -507
rect -2025 -473 -1925 -457
rect -2025 -507 -2009 -473
rect -1941 -507 -1925 -473
rect -2025 -554 -1925 -507
rect -1867 -473 -1767 -457
rect -1867 -507 -1851 -473
rect -1783 -507 -1767 -473
rect -1867 -554 -1767 -507
rect -1709 -473 -1609 -457
rect -1709 -507 -1693 -473
rect -1625 -507 -1609 -473
rect -1709 -554 -1609 -507
rect -1551 -473 -1451 -457
rect -1551 -507 -1535 -473
rect -1467 -507 -1451 -473
rect -1551 -554 -1451 -507
rect -1393 -473 -1293 -457
rect -1393 -507 -1377 -473
rect -1309 -507 -1293 -473
rect -1393 -554 -1293 -507
rect -1235 -473 -1135 -457
rect -1235 -507 -1219 -473
rect -1151 -507 -1135 -473
rect -1235 -554 -1135 -507
rect -1077 -473 -977 -457
rect -1077 -507 -1061 -473
rect -993 -507 -977 -473
rect -1077 -554 -977 -507
rect -919 -473 -819 -457
rect -919 -507 -903 -473
rect -835 -507 -819 -473
rect -919 -554 -819 -507
rect -761 -473 -661 -457
rect -761 -507 -745 -473
rect -677 -507 -661 -473
rect -761 -554 -661 -507
rect -603 -473 -503 -457
rect -603 -507 -587 -473
rect -519 -507 -503 -473
rect -603 -554 -503 -507
rect -445 -473 -345 -457
rect -445 -507 -429 -473
rect -361 -507 -345 -473
rect -445 -554 -345 -507
rect -287 -473 -187 -457
rect -287 -507 -271 -473
rect -203 -507 -187 -473
rect -287 -554 -187 -507
rect -129 -473 -29 -457
rect -129 -507 -113 -473
rect -45 -507 -29 -473
rect -129 -554 -29 -507
rect 29 -473 129 -457
rect 29 -507 45 -473
rect 113 -507 129 -473
rect 29 -554 129 -507
rect 187 -473 287 -457
rect 187 -507 203 -473
rect 271 -507 287 -473
rect 187 -554 287 -507
rect 345 -473 445 -457
rect 345 -507 361 -473
rect 429 -507 445 -473
rect 345 -554 445 -507
rect 503 -473 603 -457
rect 503 -507 519 -473
rect 587 -507 603 -473
rect 503 -554 603 -507
rect 661 -473 761 -457
rect 661 -507 677 -473
rect 745 -507 761 -473
rect 661 -554 761 -507
rect 819 -473 919 -457
rect 819 -507 835 -473
rect 903 -507 919 -473
rect 819 -554 919 -507
rect 977 -473 1077 -457
rect 977 -507 993 -473
rect 1061 -507 1077 -473
rect 977 -554 1077 -507
rect 1135 -473 1235 -457
rect 1135 -507 1151 -473
rect 1219 -507 1235 -473
rect 1135 -554 1235 -507
rect 1293 -473 1393 -457
rect 1293 -507 1309 -473
rect 1377 -507 1393 -473
rect 1293 -554 1393 -507
rect 1451 -473 1551 -457
rect 1451 -507 1467 -473
rect 1535 -507 1551 -473
rect 1451 -554 1551 -507
rect 1609 -473 1709 -457
rect 1609 -507 1625 -473
rect 1693 -507 1709 -473
rect 1609 -554 1709 -507
rect 1767 -473 1867 -457
rect 1767 -507 1783 -473
rect 1851 -507 1867 -473
rect 1767 -554 1867 -507
rect 1925 -473 2025 -457
rect 1925 -507 1941 -473
rect 2009 -507 2025 -473
rect 1925 -554 2025 -507
rect 2083 -473 2183 -457
rect 2083 -507 2099 -473
rect 2167 -507 2183 -473
rect 2083 -554 2183 -507
rect -2183 -801 -2083 -754
rect -2183 -835 -2167 -801
rect -2099 -835 -2083 -801
rect -2183 -851 -2083 -835
rect -2025 -801 -1925 -754
rect -2025 -835 -2009 -801
rect -1941 -835 -1925 -801
rect -2025 -851 -1925 -835
rect -1867 -801 -1767 -754
rect -1867 -835 -1851 -801
rect -1783 -835 -1767 -801
rect -1867 -851 -1767 -835
rect -1709 -801 -1609 -754
rect -1709 -835 -1693 -801
rect -1625 -835 -1609 -801
rect -1709 -851 -1609 -835
rect -1551 -801 -1451 -754
rect -1551 -835 -1535 -801
rect -1467 -835 -1451 -801
rect -1551 -851 -1451 -835
rect -1393 -801 -1293 -754
rect -1393 -835 -1377 -801
rect -1309 -835 -1293 -801
rect -1393 -851 -1293 -835
rect -1235 -801 -1135 -754
rect -1235 -835 -1219 -801
rect -1151 -835 -1135 -801
rect -1235 -851 -1135 -835
rect -1077 -801 -977 -754
rect -1077 -835 -1061 -801
rect -993 -835 -977 -801
rect -1077 -851 -977 -835
rect -919 -801 -819 -754
rect -919 -835 -903 -801
rect -835 -835 -819 -801
rect -919 -851 -819 -835
rect -761 -801 -661 -754
rect -761 -835 -745 -801
rect -677 -835 -661 -801
rect -761 -851 -661 -835
rect -603 -801 -503 -754
rect -603 -835 -587 -801
rect -519 -835 -503 -801
rect -603 -851 -503 -835
rect -445 -801 -345 -754
rect -445 -835 -429 -801
rect -361 -835 -345 -801
rect -445 -851 -345 -835
rect -287 -801 -187 -754
rect -287 -835 -271 -801
rect -203 -835 -187 -801
rect -287 -851 -187 -835
rect -129 -801 -29 -754
rect -129 -835 -113 -801
rect -45 -835 -29 -801
rect -129 -851 -29 -835
rect 29 -801 129 -754
rect 29 -835 45 -801
rect 113 -835 129 -801
rect 29 -851 129 -835
rect 187 -801 287 -754
rect 187 -835 203 -801
rect 271 -835 287 -801
rect 187 -851 287 -835
rect 345 -801 445 -754
rect 345 -835 361 -801
rect 429 -835 445 -801
rect 345 -851 445 -835
rect 503 -801 603 -754
rect 503 -835 519 -801
rect 587 -835 603 -801
rect 503 -851 603 -835
rect 661 -801 761 -754
rect 661 -835 677 -801
rect 745 -835 761 -801
rect 661 -851 761 -835
rect 819 -801 919 -754
rect 819 -835 835 -801
rect 903 -835 919 -801
rect 819 -851 919 -835
rect 977 -801 1077 -754
rect 977 -835 993 -801
rect 1061 -835 1077 -801
rect 977 -851 1077 -835
rect 1135 -801 1235 -754
rect 1135 -835 1151 -801
rect 1219 -835 1235 -801
rect 1135 -851 1235 -835
rect 1293 -801 1393 -754
rect 1293 -835 1309 -801
rect 1377 -835 1393 -801
rect 1293 -851 1393 -835
rect 1451 -801 1551 -754
rect 1451 -835 1467 -801
rect 1535 -835 1551 -801
rect 1451 -851 1551 -835
rect 1609 -801 1709 -754
rect 1609 -835 1625 -801
rect 1693 -835 1709 -801
rect 1609 -851 1709 -835
rect 1767 -801 1867 -754
rect 1767 -835 1783 -801
rect 1851 -835 1867 -801
rect 1767 -851 1867 -835
rect 1925 -801 2025 -754
rect 1925 -835 1941 -801
rect 2009 -835 2025 -801
rect 1925 -851 2025 -835
rect 2083 -801 2183 -754
rect 2083 -835 2099 -801
rect 2167 -835 2183 -801
rect 2083 -851 2183 -835
rect -2183 -909 -2083 -893
rect -2183 -943 -2167 -909
rect -2099 -943 -2083 -909
rect -2183 -990 -2083 -943
rect -2025 -909 -1925 -893
rect -2025 -943 -2009 -909
rect -1941 -943 -1925 -909
rect -2025 -990 -1925 -943
rect -1867 -909 -1767 -893
rect -1867 -943 -1851 -909
rect -1783 -943 -1767 -909
rect -1867 -990 -1767 -943
rect -1709 -909 -1609 -893
rect -1709 -943 -1693 -909
rect -1625 -943 -1609 -909
rect -1709 -990 -1609 -943
rect -1551 -909 -1451 -893
rect -1551 -943 -1535 -909
rect -1467 -943 -1451 -909
rect -1551 -990 -1451 -943
rect -1393 -909 -1293 -893
rect -1393 -943 -1377 -909
rect -1309 -943 -1293 -909
rect -1393 -990 -1293 -943
rect -1235 -909 -1135 -893
rect -1235 -943 -1219 -909
rect -1151 -943 -1135 -909
rect -1235 -990 -1135 -943
rect -1077 -909 -977 -893
rect -1077 -943 -1061 -909
rect -993 -943 -977 -909
rect -1077 -990 -977 -943
rect -919 -909 -819 -893
rect -919 -943 -903 -909
rect -835 -943 -819 -909
rect -919 -990 -819 -943
rect -761 -909 -661 -893
rect -761 -943 -745 -909
rect -677 -943 -661 -909
rect -761 -990 -661 -943
rect -603 -909 -503 -893
rect -603 -943 -587 -909
rect -519 -943 -503 -909
rect -603 -990 -503 -943
rect -445 -909 -345 -893
rect -445 -943 -429 -909
rect -361 -943 -345 -909
rect -445 -990 -345 -943
rect -287 -909 -187 -893
rect -287 -943 -271 -909
rect -203 -943 -187 -909
rect -287 -990 -187 -943
rect -129 -909 -29 -893
rect -129 -943 -113 -909
rect -45 -943 -29 -909
rect -129 -990 -29 -943
rect 29 -909 129 -893
rect 29 -943 45 -909
rect 113 -943 129 -909
rect 29 -990 129 -943
rect 187 -909 287 -893
rect 187 -943 203 -909
rect 271 -943 287 -909
rect 187 -990 287 -943
rect 345 -909 445 -893
rect 345 -943 361 -909
rect 429 -943 445 -909
rect 345 -990 445 -943
rect 503 -909 603 -893
rect 503 -943 519 -909
rect 587 -943 603 -909
rect 503 -990 603 -943
rect 661 -909 761 -893
rect 661 -943 677 -909
rect 745 -943 761 -909
rect 661 -990 761 -943
rect 819 -909 919 -893
rect 819 -943 835 -909
rect 903 -943 919 -909
rect 819 -990 919 -943
rect 977 -909 1077 -893
rect 977 -943 993 -909
rect 1061 -943 1077 -909
rect 977 -990 1077 -943
rect 1135 -909 1235 -893
rect 1135 -943 1151 -909
rect 1219 -943 1235 -909
rect 1135 -990 1235 -943
rect 1293 -909 1393 -893
rect 1293 -943 1309 -909
rect 1377 -943 1393 -909
rect 1293 -990 1393 -943
rect 1451 -909 1551 -893
rect 1451 -943 1467 -909
rect 1535 -943 1551 -909
rect 1451 -990 1551 -943
rect 1609 -909 1709 -893
rect 1609 -943 1625 -909
rect 1693 -943 1709 -909
rect 1609 -990 1709 -943
rect 1767 -909 1867 -893
rect 1767 -943 1783 -909
rect 1851 -943 1867 -909
rect 1767 -990 1867 -943
rect 1925 -909 2025 -893
rect 1925 -943 1941 -909
rect 2009 -943 2025 -909
rect 1925 -990 2025 -943
rect 2083 -909 2183 -893
rect 2083 -943 2099 -909
rect 2167 -943 2183 -909
rect 2083 -990 2183 -943
rect -2183 -1237 -2083 -1190
rect -2183 -1271 -2167 -1237
rect -2099 -1271 -2083 -1237
rect -2183 -1287 -2083 -1271
rect -2025 -1237 -1925 -1190
rect -2025 -1271 -2009 -1237
rect -1941 -1271 -1925 -1237
rect -2025 -1287 -1925 -1271
rect -1867 -1237 -1767 -1190
rect -1867 -1271 -1851 -1237
rect -1783 -1271 -1767 -1237
rect -1867 -1287 -1767 -1271
rect -1709 -1237 -1609 -1190
rect -1709 -1271 -1693 -1237
rect -1625 -1271 -1609 -1237
rect -1709 -1287 -1609 -1271
rect -1551 -1237 -1451 -1190
rect -1551 -1271 -1535 -1237
rect -1467 -1271 -1451 -1237
rect -1551 -1287 -1451 -1271
rect -1393 -1237 -1293 -1190
rect -1393 -1271 -1377 -1237
rect -1309 -1271 -1293 -1237
rect -1393 -1287 -1293 -1271
rect -1235 -1237 -1135 -1190
rect -1235 -1271 -1219 -1237
rect -1151 -1271 -1135 -1237
rect -1235 -1287 -1135 -1271
rect -1077 -1237 -977 -1190
rect -1077 -1271 -1061 -1237
rect -993 -1271 -977 -1237
rect -1077 -1287 -977 -1271
rect -919 -1237 -819 -1190
rect -919 -1271 -903 -1237
rect -835 -1271 -819 -1237
rect -919 -1287 -819 -1271
rect -761 -1237 -661 -1190
rect -761 -1271 -745 -1237
rect -677 -1271 -661 -1237
rect -761 -1287 -661 -1271
rect -603 -1237 -503 -1190
rect -603 -1271 -587 -1237
rect -519 -1271 -503 -1237
rect -603 -1287 -503 -1271
rect -445 -1237 -345 -1190
rect -445 -1271 -429 -1237
rect -361 -1271 -345 -1237
rect -445 -1287 -345 -1271
rect -287 -1237 -187 -1190
rect -287 -1271 -271 -1237
rect -203 -1271 -187 -1237
rect -287 -1287 -187 -1271
rect -129 -1237 -29 -1190
rect -129 -1271 -113 -1237
rect -45 -1271 -29 -1237
rect -129 -1287 -29 -1271
rect 29 -1237 129 -1190
rect 29 -1271 45 -1237
rect 113 -1271 129 -1237
rect 29 -1287 129 -1271
rect 187 -1237 287 -1190
rect 187 -1271 203 -1237
rect 271 -1271 287 -1237
rect 187 -1287 287 -1271
rect 345 -1237 445 -1190
rect 345 -1271 361 -1237
rect 429 -1271 445 -1237
rect 345 -1287 445 -1271
rect 503 -1237 603 -1190
rect 503 -1271 519 -1237
rect 587 -1271 603 -1237
rect 503 -1287 603 -1271
rect 661 -1237 761 -1190
rect 661 -1271 677 -1237
rect 745 -1271 761 -1237
rect 661 -1287 761 -1271
rect 819 -1237 919 -1190
rect 819 -1271 835 -1237
rect 903 -1271 919 -1237
rect 819 -1287 919 -1271
rect 977 -1237 1077 -1190
rect 977 -1271 993 -1237
rect 1061 -1271 1077 -1237
rect 977 -1287 1077 -1271
rect 1135 -1237 1235 -1190
rect 1135 -1271 1151 -1237
rect 1219 -1271 1235 -1237
rect 1135 -1287 1235 -1271
rect 1293 -1237 1393 -1190
rect 1293 -1271 1309 -1237
rect 1377 -1271 1393 -1237
rect 1293 -1287 1393 -1271
rect 1451 -1237 1551 -1190
rect 1451 -1271 1467 -1237
rect 1535 -1271 1551 -1237
rect 1451 -1287 1551 -1271
rect 1609 -1237 1709 -1190
rect 1609 -1271 1625 -1237
rect 1693 -1271 1709 -1237
rect 1609 -1287 1709 -1271
rect 1767 -1237 1867 -1190
rect 1767 -1271 1783 -1237
rect 1851 -1271 1867 -1237
rect 1767 -1287 1867 -1271
rect 1925 -1237 2025 -1190
rect 1925 -1271 1941 -1237
rect 2009 -1271 2025 -1237
rect 1925 -1287 2025 -1271
rect 2083 -1237 2183 -1190
rect 2083 -1271 2099 -1237
rect 2167 -1271 2183 -1237
rect 2083 -1287 2183 -1271
rect -2183 -1345 -2083 -1329
rect -2183 -1379 -2167 -1345
rect -2099 -1379 -2083 -1345
rect -2183 -1426 -2083 -1379
rect -2025 -1345 -1925 -1329
rect -2025 -1379 -2009 -1345
rect -1941 -1379 -1925 -1345
rect -2025 -1426 -1925 -1379
rect -1867 -1345 -1767 -1329
rect -1867 -1379 -1851 -1345
rect -1783 -1379 -1767 -1345
rect -1867 -1426 -1767 -1379
rect -1709 -1345 -1609 -1329
rect -1709 -1379 -1693 -1345
rect -1625 -1379 -1609 -1345
rect -1709 -1426 -1609 -1379
rect -1551 -1345 -1451 -1329
rect -1551 -1379 -1535 -1345
rect -1467 -1379 -1451 -1345
rect -1551 -1426 -1451 -1379
rect -1393 -1345 -1293 -1329
rect -1393 -1379 -1377 -1345
rect -1309 -1379 -1293 -1345
rect -1393 -1426 -1293 -1379
rect -1235 -1345 -1135 -1329
rect -1235 -1379 -1219 -1345
rect -1151 -1379 -1135 -1345
rect -1235 -1426 -1135 -1379
rect -1077 -1345 -977 -1329
rect -1077 -1379 -1061 -1345
rect -993 -1379 -977 -1345
rect -1077 -1426 -977 -1379
rect -919 -1345 -819 -1329
rect -919 -1379 -903 -1345
rect -835 -1379 -819 -1345
rect -919 -1426 -819 -1379
rect -761 -1345 -661 -1329
rect -761 -1379 -745 -1345
rect -677 -1379 -661 -1345
rect -761 -1426 -661 -1379
rect -603 -1345 -503 -1329
rect -603 -1379 -587 -1345
rect -519 -1379 -503 -1345
rect -603 -1426 -503 -1379
rect -445 -1345 -345 -1329
rect -445 -1379 -429 -1345
rect -361 -1379 -345 -1345
rect -445 -1426 -345 -1379
rect -287 -1345 -187 -1329
rect -287 -1379 -271 -1345
rect -203 -1379 -187 -1345
rect -287 -1426 -187 -1379
rect -129 -1345 -29 -1329
rect -129 -1379 -113 -1345
rect -45 -1379 -29 -1345
rect -129 -1426 -29 -1379
rect 29 -1345 129 -1329
rect 29 -1379 45 -1345
rect 113 -1379 129 -1345
rect 29 -1426 129 -1379
rect 187 -1345 287 -1329
rect 187 -1379 203 -1345
rect 271 -1379 287 -1345
rect 187 -1426 287 -1379
rect 345 -1345 445 -1329
rect 345 -1379 361 -1345
rect 429 -1379 445 -1345
rect 345 -1426 445 -1379
rect 503 -1345 603 -1329
rect 503 -1379 519 -1345
rect 587 -1379 603 -1345
rect 503 -1426 603 -1379
rect 661 -1345 761 -1329
rect 661 -1379 677 -1345
rect 745 -1379 761 -1345
rect 661 -1426 761 -1379
rect 819 -1345 919 -1329
rect 819 -1379 835 -1345
rect 903 -1379 919 -1345
rect 819 -1426 919 -1379
rect 977 -1345 1077 -1329
rect 977 -1379 993 -1345
rect 1061 -1379 1077 -1345
rect 977 -1426 1077 -1379
rect 1135 -1345 1235 -1329
rect 1135 -1379 1151 -1345
rect 1219 -1379 1235 -1345
rect 1135 -1426 1235 -1379
rect 1293 -1345 1393 -1329
rect 1293 -1379 1309 -1345
rect 1377 -1379 1393 -1345
rect 1293 -1426 1393 -1379
rect 1451 -1345 1551 -1329
rect 1451 -1379 1467 -1345
rect 1535 -1379 1551 -1345
rect 1451 -1426 1551 -1379
rect 1609 -1345 1709 -1329
rect 1609 -1379 1625 -1345
rect 1693 -1379 1709 -1345
rect 1609 -1426 1709 -1379
rect 1767 -1345 1867 -1329
rect 1767 -1379 1783 -1345
rect 1851 -1379 1867 -1345
rect 1767 -1426 1867 -1379
rect 1925 -1345 2025 -1329
rect 1925 -1379 1941 -1345
rect 2009 -1379 2025 -1345
rect 1925 -1426 2025 -1379
rect 2083 -1345 2183 -1329
rect 2083 -1379 2099 -1345
rect 2167 -1379 2183 -1345
rect 2083 -1426 2183 -1379
rect -2183 -1673 -2083 -1626
rect -2183 -1707 -2167 -1673
rect -2099 -1707 -2083 -1673
rect -2183 -1723 -2083 -1707
rect -2025 -1673 -1925 -1626
rect -2025 -1707 -2009 -1673
rect -1941 -1707 -1925 -1673
rect -2025 -1723 -1925 -1707
rect -1867 -1673 -1767 -1626
rect -1867 -1707 -1851 -1673
rect -1783 -1707 -1767 -1673
rect -1867 -1723 -1767 -1707
rect -1709 -1673 -1609 -1626
rect -1709 -1707 -1693 -1673
rect -1625 -1707 -1609 -1673
rect -1709 -1723 -1609 -1707
rect -1551 -1673 -1451 -1626
rect -1551 -1707 -1535 -1673
rect -1467 -1707 -1451 -1673
rect -1551 -1723 -1451 -1707
rect -1393 -1673 -1293 -1626
rect -1393 -1707 -1377 -1673
rect -1309 -1707 -1293 -1673
rect -1393 -1723 -1293 -1707
rect -1235 -1673 -1135 -1626
rect -1235 -1707 -1219 -1673
rect -1151 -1707 -1135 -1673
rect -1235 -1723 -1135 -1707
rect -1077 -1673 -977 -1626
rect -1077 -1707 -1061 -1673
rect -993 -1707 -977 -1673
rect -1077 -1723 -977 -1707
rect -919 -1673 -819 -1626
rect -919 -1707 -903 -1673
rect -835 -1707 -819 -1673
rect -919 -1723 -819 -1707
rect -761 -1673 -661 -1626
rect -761 -1707 -745 -1673
rect -677 -1707 -661 -1673
rect -761 -1723 -661 -1707
rect -603 -1673 -503 -1626
rect -603 -1707 -587 -1673
rect -519 -1707 -503 -1673
rect -603 -1723 -503 -1707
rect -445 -1673 -345 -1626
rect -445 -1707 -429 -1673
rect -361 -1707 -345 -1673
rect -445 -1723 -345 -1707
rect -287 -1673 -187 -1626
rect -287 -1707 -271 -1673
rect -203 -1707 -187 -1673
rect -287 -1723 -187 -1707
rect -129 -1673 -29 -1626
rect -129 -1707 -113 -1673
rect -45 -1707 -29 -1673
rect -129 -1723 -29 -1707
rect 29 -1673 129 -1626
rect 29 -1707 45 -1673
rect 113 -1707 129 -1673
rect 29 -1723 129 -1707
rect 187 -1673 287 -1626
rect 187 -1707 203 -1673
rect 271 -1707 287 -1673
rect 187 -1723 287 -1707
rect 345 -1673 445 -1626
rect 345 -1707 361 -1673
rect 429 -1707 445 -1673
rect 345 -1723 445 -1707
rect 503 -1673 603 -1626
rect 503 -1707 519 -1673
rect 587 -1707 603 -1673
rect 503 -1723 603 -1707
rect 661 -1673 761 -1626
rect 661 -1707 677 -1673
rect 745 -1707 761 -1673
rect 661 -1723 761 -1707
rect 819 -1673 919 -1626
rect 819 -1707 835 -1673
rect 903 -1707 919 -1673
rect 819 -1723 919 -1707
rect 977 -1673 1077 -1626
rect 977 -1707 993 -1673
rect 1061 -1707 1077 -1673
rect 977 -1723 1077 -1707
rect 1135 -1673 1235 -1626
rect 1135 -1707 1151 -1673
rect 1219 -1707 1235 -1673
rect 1135 -1723 1235 -1707
rect 1293 -1673 1393 -1626
rect 1293 -1707 1309 -1673
rect 1377 -1707 1393 -1673
rect 1293 -1723 1393 -1707
rect 1451 -1673 1551 -1626
rect 1451 -1707 1467 -1673
rect 1535 -1707 1551 -1673
rect 1451 -1723 1551 -1707
rect 1609 -1673 1709 -1626
rect 1609 -1707 1625 -1673
rect 1693 -1707 1709 -1673
rect 1609 -1723 1709 -1707
rect 1767 -1673 1867 -1626
rect 1767 -1707 1783 -1673
rect 1851 -1707 1867 -1673
rect 1767 -1723 1867 -1707
rect 1925 -1673 2025 -1626
rect 1925 -1707 1941 -1673
rect 2009 -1707 2025 -1673
rect 1925 -1723 2025 -1707
rect 2083 -1673 2183 -1626
rect 2083 -1707 2099 -1673
rect 2167 -1707 2183 -1673
rect 2083 -1723 2183 -1707
rect -2183 -1781 -2083 -1765
rect -2183 -1815 -2167 -1781
rect -2099 -1815 -2083 -1781
rect -2183 -1862 -2083 -1815
rect -2025 -1781 -1925 -1765
rect -2025 -1815 -2009 -1781
rect -1941 -1815 -1925 -1781
rect -2025 -1862 -1925 -1815
rect -1867 -1781 -1767 -1765
rect -1867 -1815 -1851 -1781
rect -1783 -1815 -1767 -1781
rect -1867 -1862 -1767 -1815
rect -1709 -1781 -1609 -1765
rect -1709 -1815 -1693 -1781
rect -1625 -1815 -1609 -1781
rect -1709 -1862 -1609 -1815
rect -1551 -1781 -1451 -1765
rect -1551 -1815 -1535 -1781
rect -1467 -1815 -1451 -1781
rect -1551 -1862 -1451 -1815
rect -1393 -1781 -1293 -1765
rect -1393 -1815 -1377 -1781
rect -1309 -1815 -1293 -1781
rect -1393 -1862 -1293 -1815
rect -1235 -1781 -1135 -1765
rect -1235 -1815 -1219 -1781
rect -1151 -1815 -1135 -1781
rect -1235 -1862 -1135 -1815
rect -1077 -1781 -977 -1765
rect -1077 -1815 -1061 -1781
rect -993 -1815 -977 -1781
rect -1077 -1862 -977 -1815
rect -919 -1781 -819 -1765
rect -919 -1815 -903 -1781
rect -835 -1815 -819 -1781
rect -919 -1862 -819 -1815
rect -761 -1781 -661 -1765
rect -761 -1815 -745 -1781
rect -677 -1815 -661 -1781
rect -761 -1862 -661 -1815
rect -603 -1781 -503 -1765
rect -603 -1815 -587 -1781
rect -519 -1815 -503 -1781
rect -603 -1862 -503 -1815
rect -445 -1781 -345 -1765
rect -445 -1815 -429 -1781
rect -361 -1815 -345 -1781
rect -445 -1862 -345 -1815
rect -287 -1781 -187 -1765
rect -287 -1815 -271 -1781
rect -203 -1815 -187 -1781
rect -287 -1862 -187 -1815
rect -129 -1781 -29 -1765
rect -129 -1815 -113 -1781
rect -45 -1815 -29 -1781
rect -129 -1862 -29 -1815
rect 29 -1781 129 -1765
rect 29 -1815 45 -1781
rect 113 -1815 129 -1781
rect 29 -1862 129 -1815
rect 187 -1781 287 -1765
rect 187 -1815 203 -1781
rect 271 -1815 287 -1781
rect 187 -1862 287 -1815
rect 345 -1781 445 -1765
rect 345 -1815 361 -1781
rect 429 -1815 445 -1781
rect 345 -1862 445 -1815
rect 503 -1781 603 -1765
rect 503 -1815 519 -1781
rect 587 -1815 603 -1781
rect 503 -1862 603 -1815
rect 661 -1781 761 -1765
rect 661 -1815 677 -1781
rect 745 -1815 761 -1781
rect 661 -1862 761 -1815
rect 819 -1781 919 -1765
rect 819 -1815 835 -1781
rect 903 -1815 919 -1781
rect 819 -1862 919 -1815
rect 977 -1781 1077 -1765
rect 977 -1815 993 -1781
rect 1061 -1815 1077 -1781
rect 977 -1862 1077 -1815
rect 1135 -1781 1235 -1765
rect 1135 -1815 1151 -1781
rect 1219 -1815 1235 -1781
rect 1135 -1862 1235 -1815
rect 1293 -1781 1393 -1765
rect 1293 -1815 1309 -1781
rect 1377 -1815 1393 -1781
rect 1293 -1862 1393 -1815
rect 1451 -1781 1551 -1765
rect 1451 -1815 1467 -1781
rect 1535 -1815 1551 -1781
rect 1451 -1862 1551 -1815
rect 1609 -1781 1709 -1765
rect 1609 -1815 1625 -1781
rect 1693 -1815 1709 -1781
rect 1609 -1862 1709 -1815
rect 1767 -1781 1867 -1765
rect 1767 -1815 1783 -1781
rect 1851 -1815 1867 -1781
rect 1767 -1862 1867 -1815
rect 1925 -1781 2025 -1765
rect 1925 -1815 1941 -1781
rect 2009 -1815 2025 -1781
rect 1925 -1862 2025 -1815
rect 2083 -1781 2183 -1765
rect 2083 -1815 2099 -1781
rect 2167 -1815 2183 -1781
rect 2083 -1862 2183 -1815
rect -2183 -2109 -2083 -2062
rect -2183 -2143 -2167 -2109
rect -2099 -2143 -2083 -2109
rect -2183 -2159 -2083 -2143
rect -2025 -2109 -1925 -2062
rect -2025 -2143 -2009 -2109
rect -1941 -2143 -1925 -2109
rect -2025 -2159 -1925 -2143
rect -1867 -2109 -1767 -2062
rect -1867 -2143 -1851 -2109
rect -1783 -2143 -1767 -2109
rect -1867 -2159 -1767 -2143
rect -1709 -2109 -1609 -2062
rect -1709 -2143 -1693 -2109
rect -1625 -2143 -1609 -2109
rect -1709 -2159 -1609 -2143
rect -1551 -2109 -1451 -2062
rect -1551 -2143 -1535 -2109
rect -1467 -2143 -1451 -2109
rect -1551 -2159 -1451 -2143
rect -1393 -2109 -1293 -2062
rect -1393 -2143 -1377 -2109
rect -1309 -2143 -1293 -2109
rect -1393 -2159 -1293 -2143
rect -1235 -2109 -1135 -2062
rect -1235 -2143 -1219 -2109
rect -1151 -2143 -1135 -2109
rect -1235 -2159 -1135 -2143
rect -1077 -2109 -977 -2062
rect -1077 -2143 -1061 -2109
rect -993 -2143 -977 -2109
rect -1077 -2159 -977 -2143
rect -919 -2109 -819 -2062
rect -919 -2143 -903 -2109
rect -835 -2143 -819 -2109
rect -919 -2159 -819 -2143
rect -761 -2109 -661 -2062
rect -761 -2143 -745 -2109
rect -677 -2143 -661 -2109
rect -761 -2159 -661 -2143
rect -603 -2109 -503 -2062
rect -603 -2143 -587 -2109
rect -519 -2143 -503 -2109
rect -603 -2159 -503 -2143
rect -445 -2109 -345 -2062
rect -445 -2143 -429 -2109
rect -361 -2143 -345 -2109
rect -445 -2159 -345 -2143
rect -287 -2109 -187 -2062
rect -287 -2143 -271 -2109
rect -203 -2143 -187 -2109
rect -287 -2159 -187 -2143
rect -129 -2109 -29 -2062
rect -129 -2143 -113 -2109
rect -45 -2143 -29 -2109
rect -129 -2159 -29 -2143
rect 29 -2109 129 -2062
rect 29 -2143 45 -2109
rect 113 -2143 129 -2109
rect 29 -2159 129 -2143
rect 187 -2109 287 -2062
rect 187 -2143 203 -2109
rect 271 -2143 287 -2109
rect 187 -2159 287 -2143
rect 345 -2109 445 -2062
rect 345 -2143 361 -2109
rect 429 -2143 445 -2109
rect 345 -2159 445 -2143
rect 503 -2109 603 -2062
rect 503 -2143 519 -2109
rect 587 -2143 603 -2109
rect 503 -2159 603 -2143
rect 661 -2109 761 -2062
rect 661 -2143 677 -2109
rect 745 -2143 761 -2109
rect 661 -2159 761 -2143
rect 819 -2109 919 -2062
rect 819 -2143 835 -2109
rect 903 -2143 919 -2109
rect 819 -2159 919 -2143
rect 977 -2109 1077 -2062
rect 977 -2143 993 -2109
rect 1061 -2143 1077 -2109
rect 977 -2159 1077 -2143
rect 1135 -2109 1235 -2062
rect 1135 -2143 1151 -2109
rect 1219 -2143 1235 -2109
rect 1135 -2159 1235 -2143
rect 1293 -2109 1393 -2062
rect 1293 -2143 1309 -2109
rect 1377 -2143 1393 -2109
rect 1293 -2159 1393 -2143
rect 1451 -2109 1551 -2062
rect 1451 -2143 1467 -2109
rect 1535 -2143 1551 -2109
rect 1451 -2159 1551 -2143
rect 1609 -2109 1709 -2062
rect 1609 -2143 1625 -2109
rect 1693 -2143 1709 -2109
rect 1609 -2159 1709 -2143
rect 1767 -2109 1867 -2062
rect 1767 -2143 1783 -2109
rect 1851 -2143 1867 -2109
rect 1767 -2159 1867 -2143
rect 1925 -2109 2025 -2062
rect 1925 -2143 1941 -2109
rect 2009 -2143 2025 -2109
rect 1925 -2159 2025 -2143
rect 2083 -2109 2183 -2062
rect 2083 -2143 2099 -2109
rect 2167 -2143 2183 -2109
rect 2083 -2159 2183 -2143
<< polycont >>
rect -2167 2109 -2099 2143
rect -2009 2109 -1941 2143
rect -1851 2109 -1783 2143
rect -1693 2109 -1625 2143
rect -1535 2109 -1467 2143
rect -1377 2109 -1309 2143
rect -1219 2109 -1151 2143
rect -1061 2109 -993 2143
rect -903 2109 -835 2143
rect -745 2109 -677 2143
rect -587 2109 -519 2143
rect -429 2109 -361 2143
rect -271 2109 -203 2143
rect -113 2109 -45 2143
rect 45 2109 113 2143
rect 203 2109 271 2143
rect 361 2109 429 2143
rect 519 2109 587 2143
rect 677 2109 745 2143
rect 835 2109 903 2143
rect 993 2109 1061 2143
rect 1151 2109 1219 2143
rect 1309 2109 1377 2143
rect 1467 2109 1535 2143
rect 1625 2109 1693 2143
rect 1783 2109 1851 2143
rect 1941 2109 2009 2143
rect 2099 2109 2167 2143
rect -2167 1781 -2099 1815
rect -2009 1781 -1941 1815
rect -1851 1781 -1783 1815
rect -1693 1781 -1625 1815
rect -1535 1781 -1467 1815
rect -1377 1781 -1309 1815
rect -1219 1781 -1151 1815
rect -1061 1781 -993 1815
rect -903 1781 -835 1815
rect -745 1781 -677 1815
rect -587 1781 -519 1815
rect -429 1781 -361 1815
rect -271 1781 -203 1815
rect -113 1781 -45 1815
rect 45 1781 113 1815
rect 203 1781 271 1815
rect 361 1781 429 1815
rect 519 1781 587 1815
rect 677 1781 745 1815
rect 835 1781 903 1815
rect 993 1781 1061 1815
rect 1151 1781 1219 1815
rect 1309 1781 1377 1815
rect 1467 1781 1535 1815
rect 1625 1781 1693 1815
rect 1783 1781 1851 1815
rect 1941 1781 2009 1815
rect 2099 1781 2167 1815
rect -2167 1673 -2099 1707
rect -2009 1673 -1941 1707
rect -1851 1673 -1783 1707
rect -1693 1673 -1625 1707
rect -1535 1673 -1467 1707
rect -1377 1673 -1309 1707
rect -1219 1673 -1151 1707
rect -1061 1673 -993 1707
rect -903 1673 -835 1707
rect -745 1673 -677 1707
rect -587 1673 -519 1707
rect -429 1673 -361 1707
rect -271 1673 -203 1707
rect -113 1673 -45 1707
rect 45 1673 113 1707
rect 203 1673 271 1707
rect 361 1673 429 1707
rect 519 1673 587 1707
rect 677 1673 745 1707
rect 835 1673 903 1707
rect 993 1673 1061 1707
rect 1151 1673 1219 1707
rect 1309 1673 1377 1707
rect 1467 1673 1535 1707
rect 1625 1673 1693 1707
rect 1783 1673 1851 1707
rect 1941 1673 2009 1707
rect 2099 1673 2167 1707
rect -2167 1345 -2099 1379
rect -2009 1345 -1941 1379
rect -1851 1345 -1783 1379
rect -1693 1345 -1625 1379
rect -1535 1345 -1467 1379
rect -1377 1345 -1309 1379
rect -1219 1345 -1151 1379
rect -1061 1345 -993 1379
rect -903 1345 -835 1379
rect -745 1345 -677 1379
rect -587 1345 -519 1379
rect -429 1345 -361 1379
rect -271 1345 -203 1379
rect -113 1345 -45 1379
rect 45 1345 113 1379
rect 203 1345 271 1379
rect 361 1345 429 1379
rect 519 1345 587 1379
rect 677 1345 745 1379
rect 835 1345 903 1379
rect 993 1345 1061 1379
rect 1151 1345 1219 1379
rect 1309 1345 1377 1379
rect 1467 1345 1535 1379
rect 1625 1345 1693 1379
rect 1783 1345 1851 1379
rect 1941 1345 2009 1379
rect 2099 1345 2167 1379
rect -2167 1237 -2099 1271
rect -2009 1237 -1941 1271
rect -1851 1237 -1783 1271
rect -1693 1237 -1625 1271
rect -1535 1237 -1467 1271
rect -1377 1237 -1309 1271
rect -1219 1237 -1151 1271
rect -1061 1237 -993 1271
rect -903 1237 -835 1271
rect -745 1237 -677 1271
rect -587 1237 -519 1271
rect -429 1237 -361 1271
rect -271 1237 -203 1271
rect -113 1237 -45 1271
rect 45 1237 113 1271
rect 203 1237 271 1271
rect 361 1237 429 1271
rect 519 1237 587 1271
rect 677 1237 745 1271
rect 835 1237 903 1271
rect 993 1237 1061 1271
rect 1151 1237 1219 1271
rect 1309 1237 1377 1271
rect 1467 1237 1535 1271
rect 1625 1237 1693 1271
rect 1783 1237 1851 1271
rect 1941 1237 2009 1271
rect 2099 1237 2167 1271
rect -2167 909 -2099 943
rect -2009 909 -1941 943
rect -1851 909 -1783 943
rect -1693 909 -1625 943
rect -1535 909 -1467 943
rect -1377 909 -1309 943
rect -1219 909 -1151 943
rect -1061 909 -993 943
rect -903 909 -835 943
rect -745 909 -677 943
rect -587 909 -519 943
rect -429 909 -361 943
rect -271 909 -203 943
rect -113 909 -45 943
rect 45 909 113 943
rect 203 909 271 943
rect 361 909 429 943
rect 519 909 587 943
rect 677 909 745 943
rect 835 909 903 943
rect 993 909 1061 943
rect 1151 909 1219 943
rect 1309 909 1377 943
rect 1467 909 1535 943
rect 1625 909 1693 943
rect 1783 909 1851 943
rect 1941 909 2009 943
rect 2099 909 2167 943
rect -2167 801 -2099 835
rect -2009 801 -1941 835
rect -1851 801 -1783 835
rect -1693 801 -1625 835
rect -1535 801 -1467 835
rect -1377 801 -1309 835
rect -1219 801 -1151 835
rect -1061 801 -993 835
rect -903 801 -835 835
rect -745 801 -677 835
rect -587 801 -519 835
rect -429 801 -361 835
rect -271 801 -203 835
rect -113 801 -45 835
rect 45 801 113 835
rect 203 801 271 835
rect 361 801 429 835
rect 519 801 587 835
rect 677 801 745 835
rect 835 801 903 835
rect 993 801 1061 835
rect 1151 801 1219 835
rect 1309 801 1377 835
rect 1467 801 1535 835
rect 1625 801 1693 835
rect 1783 801 1851 835
rect 1941 801 2009 835
rect 2099 801 2167 835
rect -2167 473 -2099 507
rect -2009 473 -1941 507
rect -1851 473 -1783 507
rect -1693 473 -1625 507
rect -1535 473 -1467 507
rect -1377 473 -1309 507
rect -1219 473 -1151 507
rect -1061 473 -993 507
rect -903 473 -835 507
rect -745 473 -677 507
rect -587 473 -519 507
rect -429 473 -361 507
rect -271 473 -203 507
rect -113 473 -45 507
rect 45 473 113 507
rect 203 473 271 507
rect 361 473 429 507
rect 519 473 587 507
rect 677 473 745 507
rect 835 473 903 507
rect 993 473 1061 507
rect 1151 473 1219 507
rect 1309 473 1377 507
rect 1467 473 1535 507
rect 1625 473 1693 507
rect 1783 473 1851 507
rect 1941 473 2009 507
rect 2099 473 2167 507
rect -2167 365 -2099 399
rect -2009 365 -1941 399
rect -1851 365 -1783 399
rect -1693 365 -1625 399
rect -1535 365 -1467 399
rect -1377 365 -1309 399
rect -1219 365 -1151 399
rect -1061 365 -993 399
rect -903 365 -835 399
rect -745 365 -677 399
rect -587 365 -519 399
rect -429 365 -361 399
rect -271 365 -203 399
rect -113 365 -45 399
rect 45 365 113 399
rect 203 365 271 399
rect 361 365 429 399
rect 519 365 587 399
rect 677 365 745 399
rect 835 365 903 399
rect 993 365 1061 399
rect 1151 365 1219 399
rect 1309 365 1377 399
rect 1467 365 1535 399
rect 1625 365 1693 399
rect 1783 365 1851 399
rect 1941 365 2009 399
rect 2099 365 2167 399
rect -2167 37 -2099 71
rect -2009 37 -1941 71
rect -1851 37 -1783 71
rect -1693 37 -1625 71
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect 1625 37 1693 71
rect 1783 37 1851 71
rect 1941 37 2009 71
rect 2099 37 2167 71
rect -2167 -71 -2099 -37
rect -2009 -71 -1941 -37
rect -1851 -71 -1783 -37
rect -1693 -71 -1625 -37
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect 1625 -71 1693 -37
rect 1783 -71 1851 -37
rect 1941 -71 2009 -37
rect 2099 -71 2167 -37
rect -2167 -399 -2099 -365
rect -2009 -399 -1941 -365
rect -1851 -399 -1783 -365
rect -1693 -399 -1625 -365
rect -1535 -399 -1467 -365
rect -1377 -399 -1309 -365
rect -1219 -399 -1151 -365
rect -1061 -399 -993 -365
rect -903 -399 -835 -365
rect -745 -399 -677 -365
rect -587 -399 -519 -365
rect -429 -399 -361 -365
rect -271 -399 -203 -365
rect -113 -399 -45 -365
rect 45 -399 113 -365
rect 203 -399 271 -365
rect 361 -399 429 -365
rect 519 -399 587 -365
rect 677 -399 745 -365
rect 835 -399 903 -365
rect 993 -399 1061 -365
rect 1151 -399 1219 -365
rect 1309 -399 1377 -365
rect 1467 -399 1535 -365
rect 1625 -399 1693 -365
rect 1783 -399 1851 -365
rect 1941 -399 2009 -365
rect 2099 -399 2167 -365
rect -2167 -507 -2099 -473
rect -2009 -507 -1941 -473
rect -1851 -507 -1783 -473
rect -1693 -507 -1625 -473
rect -1535 -507 -1467 -473
rect -1377 -507 -1309 -473
rect -1219 -507 -1151 -473
rect -1061 -507 -993 -473
rect -903 -507 -835 -473
rect -745 -507 -677 -473
rect -587 -507 -519 -473
rect -429 -507 -361 -473
rect -271 -507 -203 -473
rect -113 -507 -45 -473
rect 45 -507 113 -473
rect 203 -507 271 -473
rect 361 -507 429 -473
rect 519 -507 587 -473
rect 677 -507 745 -473
rect 835 -507 903 -473
rect 993 -507 1061 -473
rect 1151 -507 1219 -473
rect 1309 -507 1377 -473
rect 1467 -507 1535 -473
rect 1625 -507 1693 -473
rect 1783 -507 1851 -473
rect 1941 -507 2009 -473
rect 2099 -507 2167 -473
rect -2167 -835 -2099 -801
rect -2009 -835 -1941 -801
rect -1851 -835 -1783 -801
rect -1693 -835 -1625 -801
rect -1535 -835 -1467 -801
rect -1377 -835 -1309 -801
rect -1219 -835 -1151 -801
rect -1061 -835 -993 -801
rect -903 -835 -835 -801
rect -745 -835 -677 -801
rect -587 -835 -519 -801
rect -429 -835 -361 -801
rect -271 -835 -203 -801
rect -113 -835 -45 -801
rect 45 -835 113 -801
rect 203 -835 271 -801
rect 361 -835 429 -801
rect 519 -835 587 -801
rect 677 -835 745 -801
rect 835 -835 903 -801
rect 993 -835 1061 -801
rect 1151 -835 1219 -801
rect 1309 -835 1377 -801
rect 1467 -835 1535 -801
rect 1625 -835 1693 -801
rect 1783 -835 1851 -801
rect 1941 -835 2009 -801
rect 2099 -835 2167 -801
rect -2167 -943 -2099 -909
rect -2009 -943 -1941 -909
rect -1851 -943 -1783 -909
rect -1693 -943 -1625 -909
rect -1535 -943 -1467 -909
rect -1377 -943 -1309 -909
rect -1219 -943 -1151 -909
rect -1061 -943 -993 -909
rect -903 -943 -835 -909
rect -745 -943 -677 -909
rect -587 -943 -519 -909
rect -429 -943 -361 -909
rect -271 -943 -203 -909
rect -113 -943 -45 -909
rect 45 -943 113 -909
rect 203 -943 271 -909
rect 361 -943 429 -909
rect 519 -943 587 -909
rect 677 -943 745 -909
rect 835 -943 903 -909
rect 993 -943 1061 -909
rect 1151 -943 1219 -909
rect 1309 -943 1377 -909
rect 1467 -943 1535 -909
rect 1625 -943 1693 -909
rect 1783 -943 1851 -909
rect 1941 -943 2009 -909
rect 2099 -943 2167 -909
rect -2167 -1271 -2099 -1237
rect -2009 -1271 -1941 -1237
rect -1851 -1271 -1783 -1237
rect -1693 -1271 -1625 -1237
rect -1535 -1271 -1467 -1237
rect -1377 -1271 -1309 -1237
rect -1219 -1271 -1151 -1237
rect -1061 -1271 -993 -1237
rect -903 -1271 -835 -1237
rect -745 -1271 -677 -1237
rect -587 -1271 -519 -1237
rect -429 -1271 -361 -1237
rect -271 -1271 -203 -1237
rect -113 -1271 -45 -1237
rect 45 -1271 113 -1237
rect 203 -1271 271 -1237
rect 361 -1271 429 -1237
rect 519 -1271 587 -1237
rect 677 -1271 745 -1237
rect 835 -1271 903 -1237
rect 993 -1271 1061 -1237
rect 1151 -1271 1219 -1237
rect 1309 -1271 1377 -1237
rect 1467 -1271 1535 -1237
rect 1625 -1271 1693 -1237
rect 1783 -1271 1851 -1237
rect 1941 -1271 2009 -1237
rect 2099 -1271 2167 -1237
rect -2167 -1379 -2099 -1345
rect -2009 -1379 -1941 -1345
rect -1851 -1379 -1783 -1345
rect -1693 -1379 -1625 -1345
rect -1535 -1379 -1467 -1345
rect -1377 -1379 -1309 -1345
rect -1219 -1379 -1151 -1345
rect -1061 -1379 -993 -1345
rect -903 -1379 -835 -1345
rect -745 -1379 -677 -1345
rect -587 -1379 -519 -1345
rect -429 -1379 -361 -1345
rect -271 -1379 -203 -1345
rect -113 -1379 -45 -1345
rect 45 -1379 113 -1345
rect 203 -1379 271 -1345
rect 361 -1379 429 -1345
rect 519 -1379 587 -1345
rect 677 -1379 745 -1345
rect 835 -1379 903 -1345
rect 993 -1379 1061 -1345
rect 1151 -1379 1219 -1345
rect 1309 -1379 1377 -1345
rect 1467 -1379 1535 -1345
rect 1625 -1379 1693 -1345
rect 1783 -1379 1851 -1345
rect 1941 -1379 2009 -1345
rect 2099 -1379 2167 -1345
rect -2167 -1707 -2099 -1673
rect -2009 -1707 -1941 -1673
rect -1851 -1707 -1783 -1673
rect -1693 -1707 -1625 -1673
rect -1535 -1707 -1467 -1673
rect -1377 -1707 -1309 -1673
rect -1219 -1707 -1151 -1673
rect -1061 -1707 -993 -1673
rect -903 -1707 -835 -1673
rect -745 -1707 -677 -1673
rect -587 -1707 -519 -1673
rect -429 -1707 -361 -1673
rect -271 -1707 -203 -1673
rect -113 -1707 -45 -1673
rect 45 -1707 113 -1673
rect 203 -1707 271 -1673
rect 361 -1707 429 -1673
rect 519 -1707 587 -1673
rect 677 -1707 745 -1673
rect 835 -1707 903 -1673
rect 993 -1707 1061 -1673
rect 1151 -1707 1219 -1673
rect 1309 -1707 1377 -1673
rect 1467 -1707 1535 -1673
rect 1625 -1707 1693 -1673
rect 1783 -1707 1851 -1673
rect 1941 -1707 2009 -1673
rect 2099 -1707 2167 -1673
rect -2167 -1815 -2099 -1781
rect -2009 -1815 -1941 -1781
rect -1851 -1815 -1783 -1781
rect -1693 -1815 -1625 -1781
rect -1535 -1815 -1467 -1781
rect -1377 -1815 -1309 -1781
rect -1219 -1815 -1151 -1781
rect -1061 -1815 -993 -1781
rect -903 -1815 -835 -1781
rect -745 -1815 -677 -1781
rect -587 -1815 -519 -1781
rect -429 -1815 -361 -1781
rect -271 -1815 -203 -1781
rect -113 -1815 -45 -1781
rect 45 -1815 113 -1781
rect 203 -1815 271 -1781
rect 361 -1815 429 -1781
rect 519 -1815 587 -1781
rect 677 -1815 745 -1781
rect 835 -1815 903 -1781
rect 993 -1815 1061 -1781
rect 1151 -1815 1219 -1781
rect 1309 -1815 1377 -1781
rect 1467 -1815 1535 -1781
rect 1625 -1815 1693 -1781
rect 1783 -1815 1851 -1781
rect 1941 -1815 2009 -1781
rect 2099 -1815 2167 -1781
rect -2167 -2143 -2099 -2109
rect -2009 -2143 -1941 -2109
rect -1851 -2143 -1783 -2109
rect -1693 -2143 -1625 -2109
rect -1535 -2143 -1467 -2109
rect -1377 -2143 -1309 -2109
rect -1219 -2143 -1151 -2109
rect -1061 -2143 -993 -2109
rect -903 -2143 -835 -2109
rect -745 -2143 -677 -2109
rect -587 -2143 -519 -2109
rect -429 -2143 -361 -2109
rect -271 -2143 -203 -2109
rect -113 -2143 -45 -2109
rect 45 -2143 113 -2109
rect 203 -2143 271 -2109
rect 361 -2143 429 -2109
rect 519 -2143 587 -2109
rect 677 -2143 745 -2109
rect 835 -2143 903 -2109
rect 993 -2143 1061 -2109
rect 1151 -2143 1219 -2109
rect 1309 -2143 1377 -2109
rect 1467 -2143 1535 -2109
rect 1625 -2143 1693 -2109
rect 1783 -2143 1851 -2109
rect 1941 -2143 2009 -2109
rect 2099 -2143 2167 -2109
<< locali >>
rect -2363 2247 -2267 2281
rect 2267 2247 2363 2281
rect -2363 2185 -2329 2247
rect 2329 2185 2363 2247
rect -2183 2109 -2167 2143
rect -2099 2109 -2083 2143
rect -2025 2109 -2009 2143
rect -1941 2109 -1925 2143
rect -1867 2109 -1851 2143
rect -1783 2109 -1767 2143
rect -1709 2109 -1693 2143
rect -1625 2109 -1609 2143
rect -1551 2109 -1535 2143
rect -1467 2109 -1451 2143
rect -1393 2109 -1377 2143
rect -1309 2109 -1293 2143
rect -1235 2109 -1219 2143
rect -1151 2109 -1135 2143
rect -1077 2109 -1061 2143
rect -993 2109 -977 2143
rect -919 2109 -903 2143
rect -835 2109 -819 2143
rect -761 2109 -745 2143
rect -677 2109 -661 2143
rect -603 2109 -587 2143
rect -519 2109 -503 2143
rect -445 2109 -429 2143
rect -361 2109 -345 2143
rect -287 2109 -271 2143
rect -203 2109 -187 2143
rect -129 2109 -113 2143
rect -45 2109 -29 2143
rect 29 2109 45 2143
rect 113 2109 129 2143
rect 187 2109 203 2143
rect 271 2109 287 2143
rect 345 2109 361 2143
rect 429 2109 445 2143
rect 503 2109 519 2143
rect 587 2109 603 2143
rect 661 2109 677 2143
rect 745 2109 761 2143
rect 819 2109 835 2143
rect 903 2109 919 2143
rect 977 2109 993 2143
rect 1061 2109 1077 2143
rect 1135 2109 1151 2143
rect 1219 2109 1235 2143
rect 1293 2109 1309 2143
rect 1377 2109 1393 2143
rect 1451 2109 1467 2143
rect 1535 2109 1551 2143
rect 1609 2109 1625 2143
rect 1693 2109 1709 2143
rect 1767 2109 1783 2143
rect 1851 2109 1867 2143
rect 1925 2109 1941 2143
rect 2009 2109 2025 2143
rect 2083 2109 2099 2143
rect 2167 2109 2183 2143
rect -2229 2050 -2195 2066
rect -2229 1858 -2195 1874
rect -2071 2050 -2037 2066
rect -2071 1858 -2037 1874
rect -1913 2050 -1879 2066
rect -1913 1858 -1879 1874
rect -1755 2050 -1721 2066
rect -1755 1858 -1721 1874
rect -1597 2050 -1563 2066
rect -1597 1858 -1563 1874
rect -1439 2050 -1405 2066
rect -1439 1858 -1405 1874
rect -1281 2050 -1247 2066
rect -1281 1858 -1247 1874
rect -1123 2050 -1089 2066
rect -1123 1858 -1089 1874
rect -965 2050 -931 2066
rect -965 1858 -931 1874
rect -807 2050 -773 2066
rect -807 1858 -773 1874
rect -649 2050 -615 2066
rect -649 1858 -615 1874
rect -491 2050 -457 2066
rect -491 1858 -457 1874
rect -333 2050 -299 2066
rect -333 1858 -299 1874
rect -175 2050 -141 2066
rect -175 1858 -141 1874
rect -17 2050 17 2066
rect -17 1858 17 1874
rect 141 2050 175 2066
rect 141 1858 175 1874
rect 299 2050 333 2066
rect 299 1858 333 1874
rect 457 2050 491 2066
rect 457 1858 491 1874
rect 615 2050 649 2066
rect 615 1858 649 1874
rect 773 2050 807 2066
rect 773 1858 807 1874
rect 931 2050 965 2066
rect 931 1858 965 1874
rect 1089 2050 1123 2066
rect 1089 1858 1123 1874
rect 1247 2050 1281 2066
rect 1247 1858 1281 1874
rect 1405 2050 1439 2066
rect 1405 1858 1439 1874
rect 1563 2050 1597 2066
rect 1563 1858 1597 1874
rect 1721 2050 1755 2066
rect 1721 1858 1755 1874
rect 1879 2050 1913 2066
rect 1879 1858 1913 1874
rect 2037 2050 2071 2066
rect 2037 1858 2071 1874
rect 2195 2050 2229 2066
rect 2195 1858 2229 1874
rect -2183 1781 -2167 1815
rect -2099 1781 -2083 1815
rect -2025 1781 -2009 1815
rect -1941 1781 -1925 1815
rect -1867 1781 -1851 1815
rect -1783 1781 -1767 1815
rect -1709 1781 -1693 1815
rect -1625 1781 -1609 1815
rect -1551 1781 -1535 1815
rect -1467 1781 -1451 1815
rect -1393 1781 -1377 1815
rect -1309 1781 -1293 1815
rect -1235 1781 -1219 1815
rect -1151 1781 -1135 1815
rect -1077 1781 -1061 1815
rect -993 1781 -977 1815
rect -919 1781 -903 1815
rect -835 1781 -819 1815
rect -761 1781 -745 1815
rect -677 1781 -661 1815
rect -603 1781 -587 1815
rect -519 1781 -503 1815
rect -445 1781 -429 1815
rect -361 1781 -345 1815
rect -287 1781 -271 1815
rect -203 1781 -187 1815
rect -129 1781 -113 1815
rect -45 1781 -29 1815
rect 29 1781 45 1815
rect 113 1781 129 1815
rect 187 1781 203 1815
rect 271 1781 287 1815
rect 345 1781 361 1815
rect 429 1781 445 1815
rect 503 1781 519 1815
rect 587 1781 603 1815
rect 661 1781 677 1815
rect 745 1781 761 1815
rect 819 1781 835 1815
rect 903 1781 919 1815
rect 977 1781 993 1815
rect 1061 1781 1077 1815
rect 1135 1781 1151 1815
rect 1219 1781 1235 1815
rect 1293 1781 1309 1815
rect 1377 1781 1393 1815
rect 1451 1781 1467 1815
rect 1535 1781 1551 1815
rect 1609 1781 1625 1815
rect 1693 1781 1709 1815
rect 1767 1781 1783 1815
rect 1851 1781 1867 1815
rect 1925 1781 1941 1815
rect 2009 1781 2025 1815
rect 2083 1781 2099 1815
rect 2167 1781 2183 1815
rect -2183 1673 -2167 1707
rect -2099 1673 -2083 1707
rect -2025 1673 -2009 1707
rect -1941 1673 -1925 1707
rect -1867 1673 -1851 1707
rect -1783 1673 -1767 1707
rect -1709 1673 -1693 1707
rect -1625 1673 -1609 1707
rect -1551 1673 -1535 1707
rect -1467 1673 -1451 1707
rect -1393 1673 -1377 1707
rect -1309 1673 -1293 1707
rect -1235 1673 -1219 1707
rect -1151 1673 -1135 1707
rect -1077 1673 -1061 1707
rect -993 1673 -977 1707
rect -919 1673 -903 1707
rect -835 1673 -819 1707
rect -761 1673 -745 1707
rect -677 1673 -661 1707
rect -603 1673 -587 1707
rect -519 1673 -503 1707
rect -445 1673 -429 1707
rect -361 1673 -345 1707
rect -287 1673 -271 1707
rect -203 1673 -187 1707
rect -129 1673 -113 1707
rect -45 1673 -29 1707
rect 29 1673 45 1707
rect 113 1673 129 1707
rect 187 1673 203 1707
rect 271 1673 287 1707
rect 345 1673 361 1707
rect 429 1673 445 1707
rect 503 1673 519 1707
rect 587 1673 603 1707
rect 661 1673 677 1707
rect 745 1673 761 1707
rect 819 1673 835 1707
rect 903 1673 919 1707
rect 977 1673 993 1707
rect 1061 1673 1077 1707
rect 1135 1673 1151 1707
rect 1219 1673 1235 1707
rect 1293 1673 1309 1707
rect 1377 1673 1393 1707
rect 1451 1673 1467 1707
rect 1535 1673 1551 1707
rect 1609 1673 1625 1707
rect 1693 1673 1709 1707
rect 1767 1673 1783 1707
rect 1851 1673 1867 1707
rect 1925 1673 1941 1707
rect 2009 1673 2025 1707
rect 2083 1673 2099 1707
rect 2167 1673 2183 1707
rect -2229 1614 -2195 1630
rect -2229 1422 -2195 1438
rect -2071 1614 -2037 1630
rect -2071 1422 -2037 1438
rect -1913 1614 -1879 1630
rect -1913 1422 -1879 1438
rect -1755 1614 -1721 1630
rect -1755 1422 -1721 1438
rect -1597 1614 -1563 1630
rect -1597 1422 -1563 1438
rect -1439 1614 -1405 1630
rect -1439 1422 -1405 1438
rect -1281 1614 -1247 1630
rect -1281 1422 -1247 1438
rect -1123 1614 -1089 1630
rect -1123 1422 -1089 1438
rect -965 1614 -931 1630
rect -965 1422 -931 1438
rect -807 1614 -773 1630
rect -807 1422 -773 1438
rect -649 1614 -615 1630
rect -649 1422 -615 1438
rect -491 1614 -457 1630
rect -491 1422 -457 1438
rect -333 1614 -299 1630
rect -333 1422 -299 1438
rect -175 1614 -141 1630
rect -175 1422 -141 1438
rect -17 1614 17 1630
rect -17 1422 17 1438
rect 141 1614 175 1630
rect 141 1422 175 1438
rect 299 1614 333 1630
rect 299 1422 333 1438
rect 457 1614 491 1630
rect 457 1422 491 1438
rect 615 1614 649 1630
rect 615 1422 649 1438
rect 773 1614 807 1630
rect 773 1422 807 1438
rect 931 1614 965 1630
rect 931 1422 965 1438
rect 1089 1614 1123 1630
rect 1089 1422 1123 1438
rect 1247 1614 1281 1630
rect 1247 1422 1281 1438
rect 1405 1614 1439 1630
rect 1405 1422 1439 1438
rect 1563 1614 1597 1630
rect 1563 1422 1597 1438
rect 1721 1614 1755 1630
rect 1721 1422 1755 1438
rect 1879 1614 1913 1630
rect 1879 1422 1913 1438
rect 2037 1614 2071 1630
rect 2037 1422 2071 1438
rect 2195 1614 2229 1630
rect 2195 1422 2229 1438
rect -2183 1345 -2167 1379
rect -2099 1345 -2083 1379
rect -2025 1345 -2009 1379
rect -1941 1345 -1925 1379
rect -1867 1345 -1851 1379
rect -1783 1345 -1767 1379
rect -1709 1345 -1693 1379
rect -1625 1345 -1609 1379
rect -1551 1345 -1535 1379
rect -1467 1345 -1451 1379
rect -1393 1345 -1377 1379
rect -1309 1345 -1293 1379
rect -1235 1345 -1219 1379
rect -1151 1345 -1135 1379
rect -1077 1345 -1061 1379
rect -993 1345 -977 1379
rect -919 1345 -903 1379
rect -835 1345 -819 1379
rect -761 1345 -745 1379
rect -677 1345 -661 1379
rect -603 1345 -587 1379
rect -519 1345 -503 1379
rect -445 1345 -429 1379
rect -361 1345 -345 1379
rect -287 1345 -271 1379
rect -203 1345 -187 1379
rect -129 1345 -113 1379
rect -45 1345 -29 1379
rect 29 1345 45 1379
rect 113 1345 129 1379
rect 187 1345 203 1379
rect 271 1345 287 1379
rect 345 1345 361 1379
rect 429 1345 445 1379
rect 503 1345 519 1379
rect 587 1345 603 1379
rect 661 1345 677 1379
rect 745 1345 761 1379
rect 819 1345 835 1379
rect 903 1345 919 1379
rect 977 1345 993 1379
rect 1061 1345 1077 1379
rect 1135 1345 1151 1379
rect 1219 1345 1235 1379
rect 1293 1345 1309 1379
rect 1377 1345 1393 1379
rect 1451 1345 1467 1379
rect 1535 1345 1551 1379
rect 1609 1345 1625 1379
rect 1693 1345 1709 1379
rect 1767 1345 1783 1379
rect 1851 1345 1867 1379
rect 1925 1345 1941 1379
rect 2009 1345 2025 1379
rect 2083 1345 2099 1379
rect 2167 1345 2183 1379
rect -2183 1237 -2167 1271
rect -2099 1237 -2083 1271
rect -2025 1237 -2009 1271
rect -1941 1237 -1925 1271
rect -1867 1237 -1851 1271
rect -1783 1237 -1767 1271
rect -1709 1237 -1693 1271
rect -1625 1237 -1609 1271
rect -1551 1237 -1535 1271
rect -1467 1237 -1451 1271
rect -1393 1237 -1377 1271
rect -1309 1237 -1293 1271
rect -1235 1237 -1219 1271
rect -1151 1237 -1135 1271
rect -1077 1237 -1061 1271
rect -993 1237 -977 1271
rect -919 1237 -903 1271
rect -835 1237 -819 1271
rect -761 1237 -745 1271
rect -677 1237 -661 1271
rect -603 1237 -587 1271
rect -519 1237 -503 1271
rect -445 1237 -429 1271
rect -361 1237 -345 1271
rect -287 1237 -271 1271
rect -203 1237 -187 1271
rect -129 1237 -113 1271
rect -45 1237 -29 1271
rect 29 1237 45 1271
rect 113 1237 129 1271
rect 187 1237 203 1271
rect 271 1237 287 1271
rect 345 1237 361 1271
rect 429 1237 445 1271
rect 503 1237 519 1271
rect 587 1237 603 1271
rect 661 1237 677 1271
rect 745 1237 761 1271
rect 819 1237 835 1271
rect 903 1237 919 1271
rect 977 1237 993 1271
rect 1061 1237 1077 1271
rect 1135 1237 1151 1271
rect 1219 1237 1235 1271
rect 1293 1237 1309 1271
rect 1377 1237 1393 1271
rect 1451 1237 1467 1271
rect 1535 1237 1551 1271
rect 1609 1237 1625 1271
rect 1693 1237 1709 1271
rect 1767 1237 1783 1271
rect 1851 1237 1867 1271
rect 1925 1237 1941 1271
rect 2009 1237 2025 1271
rect 2083 1237 2099 1271
rect 2167 1237 2183 1271
rect -2229 1178 -2195 1194
rect -2229 986 -2195 1002
rect -2071 1178 -2037 1194
rect -2071 986 -2037 1002
rect -1913 1178 -1879 1194
rect -1913 986 -1879 1002
rect -1755 1178 -1721 1194
rect -1755 986 -1721 1002
rect -1597 1178 -1563 1194
rect -1597 986 -1563 1002
rect -1439 1178 -1405 1194
rect -1439 986 -1405 1002
rect -1281 1178 -1247 1194
rect -1281 986 -1247 1002
rect -1123 1178 -1089 1194
rect -1123 986 -1089 1002
rect -965 1178 -931 1194
rect -965 986 -931 1002
rect -807 1178 -773 1194
rect -807 986 -773 1002
rect -649 1178 -615 1194
rect -649 986 -615 1002
rect -491 1178 -457 1194
rect -491 986 -457 1002
rect -333 1178 -299 1194
rect -333 986 -299 1002
rect -175 1178 -141 1194
rect -175 986 -141 1002
rect -17 1178 17 1194
rect -17 986 17 1002
rect 141 1178 175 1194
rect 141 986 175 1002
rect 299 1178 333 1194
rect 299 986 333 1002
rect 457 1178 491 1194
rect 457 986 491 1002
rect 615 1178 649 1194
rect 615 986 649 1002
rect 773 1178 807 1194
rect 773 986 807 1002
rect 931 1178 965 1194
rect 931 986 965 1002
rect 1089 1178 1123 1194
rect 1089 986 1123 1002
rect 1247 1178 1281 1194
rect 1247 986 1281 1002
rect 1405 1178 1439 1194
rect 1405 986 1439 1002
rect 1563 1178 1597 1194
rect 1563 986 1597 1002
rect 1721 1178 1755 1194
rect 1721 986 1755 1002
rect 1879 1178 1913 1194
rect 1879 986 1913 1002
rect 2037 1178 2071 1194
rect 2037 986 2071 1002
rect 2195 1178 2229 1194
rect 2195 986 2229 1002
rect -2183 909 -2167 943
rect -2099 909 -2083 943
rect -2025 909 -2009 943
rect -1941 909 -1925 943
rect -1867 909 -1851 943
rect -1783 909 -1767 943
rect -1709 909 -1693 943
rect -1625 909 -1609 943
rect -1551 909 -1535 943
rect -1467 909 -1451 943
rect -1393 909 -1377 943
rect -1309 909 -1293 943
rect -1235 909 -1219 943
rect -1151 909 -1135 943
rect -1077 909 -1061 943
rect -993 909 -977 943
rect -919 909 -903 943
rect -835 909 -819 943
rect -761 909 -745 943
rect -677 909 -661 943
rect -603 909 -587 943
rect -519 909 -503 943
rect -445 909 -429 943
rect -361 909 -345 943
rect -287 909 -271 943
rect -203 909 -187 943
rect -129 909 -113 943
rect -45 909 -29 943
rect 29 909 45 943
rect 113 909 129 943
rect 187 909 203 943
rect 271 909 287 943
rect 345 909 361 943
rect 429 909 445 943
rect 503 909 519 943
rect 587 909 603 943
rect 661 909 677 943
rect 745 909 761 943
rect 819 909 835 943
rect 903 909 919 943
rect 977 909 993 943
rect 1061 909 1077 943
rect 1135 909 1151 943
rect 1219 909 1235 943
rect 1293 909 1309 943
rect 1377 909 1393 943
rect 1451 909 1467 943
rect 1535 909 1551 943
rect 1609 909 1625 943
rect 1693 909 1709 943
rect 1767 909 1783 943
rect 1851 909 1867 943
rect 1925 909 1941 943
rect 2009 909 2025 943
rect 2083 909 2099 943
rect 2167 909 2183 943
rect -2183 801 -2167 835
rect -2099 801 -2083 835
rect -2025 801 -2009 835
rect -1941 801 -1925 835
rect -1867 801 -1851 835
rect -1783 801 -1767 835
rect -1709 801 -1693 835
rect -1625 801 -1609 835
rect -1551 801 -1535 835
rect -1467 801 -1451 835
rect -1393 801 -1377 835
rect -1309 801 -1293 835
rect -1235 801 -1219 835
rect -1151 801 -1135 835
rect -1077 801 -1061 835
rect -993 801 -977 835
rect -919 801 -903 835
rect -835 801 -819 835
rect -761 801 -745 835
rect -677 801 -661 835
rect -603 801 -587 835
rect -519 801 -503 835
rect -445 801 -429 835
rect -361 801 -345 835
rect -287 801 -271 835
rect -203 801 -187 835
rect -129 801 -113 835
rect -45 801 -29 835
rect 29 801 45 835
rect 113 801 129 835
rect 187 801 203 835
rect 271 801 287 835
rect 345 801 361 835
rect 429 801 445 835
rect 503 801 519 835
rect 587 801 603 835
rect 661 801 677 835
rect 745 801 761 835
rect 819 801 835 835
rect 903 801 919 835
rect 977 801 993 835
rect 1061 801 1077 835
rect 1135 801 1151 835
rect 1219 801 1235 835
rect 1293 801 1309 835
rect 1377 801 1393 835
rect 1451 801 1467 835
rect 1535 801 1551 835
rect 1609 801 1625 835
rect 1693 801 1709 835
rect 1767 801 1783 835
rect 1851 801 1867 835
rect 1925 801 1941 835
rect 2009 801 2025 835
rect 2083 801 2099 835
rect 2167 801 2183 835
rect -2229 742 -2195 758
rect -2229 550 -2195 566
rect -2071 742 -2037 758
rect -2071 550 -2037 566
rect -1913 742 -1879 758
rect -1913 550 -1879 566
rect -1755 742 -1721 758
rect -1755 550 -1721 566
rect -1597 742 -1563 758
rect -1597 550 -1563 566
rect -1439 742 -1405 758
rect -1439 550 -1405 566
rect -1281 742 -1247 758
rect -1281 550 -1247 566
rect -1123 742 -1089 758
rect -1123 550 -1089 566
rect -965 742 -931 758
rect -965 550 -931 566
rect -807 742 -773 758
rect -807 550 -773 566
rect -649 742 -615 758
rect -649 550 -615 566
rect -491 742 -457 758
rect -491 550 -457 566
rect -333 742 -299 758
rect -333 550 -299 566
rect -175 742 -141 758
rect -175 550 -141 566
rect -17 742 17 758
rect -17 550 17 566
rect 141 742 175 758
rect 141 550 175 566
rect 299 742 333 758
rect 299 550 333 566
rect 457 742 491 758
rect 457 550 491 566
rect 615 742 649 758
rect 615 550 649 566
rect 773 742 807 758
rect 773 550 807 566
rect 931 742 965 758
rect 931 550 965 566
rect 1089 742 1123 758
rect 1089 550 1123 566
rect 1247 742 1281 758
rect 1247 550 1281 566
rect 1405 742 1439 758
rect 1405 550 1439 566
rect 1563 742 1597 758
rect 1563 550 1597 566
rect 1721 742 1755 758
rect 1721 550 1755 566
rect 1879 742 1913 758
rect 1879 550 1913 566
rect 2037 742 2071 758
rect 2037 550 2071 566
rect 2195 742 2229 758
rect 2195 550 2229 566
rect -2183 473 -2167 507
rect -2099 473 -2083 507
rect -2025 473 -2009 507
rect -1941 473 -1925 507
rect -1867 473 -1851 507
rect -1783 473 -1767 507
rect -1709 473 -1693 507
rect -1625 473 -1609 507
rect -1551 473 -1535 507
rect -1467 473 -1451 507
rect -1393 473 -1377 507
rect -1309 473 -1293 507
rect -1235 473 -1219 507
rect -1151 473 -1135 507
rect -1077 473 -1061 507
rect -993 473 -977 507
rect -919 473 -903 507
rect -835 473 -819 507
rect -761 473 -745 507
rect -677 473 -661 507
rect -603 473 -587 507
rect -519 473 -503 507
rect -445 473 -429 507
rect -361 473 -345 507
rect -287 473 -271 507
rect -203 473 -187 507
rect -129 473 -113 507
rect -45 473 -29 507
rect 29 473 45 507
rect 113 473 129 507
rect 187 473 203 507
rect 271 473 287 507
rect 345 473 361 507
rect 429 473 445 507
rect 503 473 519 507
rect 587 473 603 507
rect 661 473 677 507
rect 745 473 761 507
rect 819 473 835 507
rect 903 473 919 507
rect 977 473 993 507
rect 1061 473 1077 507
rect 1135 473 1151 507
rect 1219 473 1235 507
rect 1293 473 1309 507
rect 1377 473 1393 507
rect 1451 473 1467 507
rect 1535 473 1551 507
rect 1609 473 1625 507
rect 1693 473 1709 507
rect 1767 473 1783 507
rect 1851 473 1867 507
rect 1925 473 1941 507
rect 2009 473 2025 507
rect 2083 473 2099 507
rect 2167 473 2183 507
rect -2183 365 -2167 399
rect -2099 365 -2083 399
rect -2025 365 -2009 399
rect -1941 365 -1925 399
rect -1867 365 -1851 399
rect -1783 365 -1767 399
rect -1709 365 -1693 399
rect -1625 365 -1609 399
rect -1551 365 -1535 399
rect -1467 365 -1451 399
rect -1393 365 -1377 399
rect -1309 365 -1293 399
rect -1235 365 -1219 399
rect -1151 365 -1135 399
rect -1077 365 -1061 399
rect -993 365 -977 399
rect -919 365 -903 399
rect -835 365 -819 399
rect -761 365 -745 399
rect -677 365 -661 399
rect -603 365 -587 399
rect -519 365 -503 399
rect -445 365 -429 399
rect -361 365 -345 399
rect -287 365 -271 399
rect -203 365 -187 399
rect -129 365 -113 399
rect -45 365 -29 399
rect 29 365 45 399
rect 113 365 129 399
rect 187 365 203 399
rect 271 365 287 399
rect 345 365 361 399
rect 429 365 445 399
rect 503 365 519 399
rect 587 365 603 399
rect 661 365 677 399
rect 745 365 761 399
rect 819 365 835 399
rect 903 365 919 399
rect 977 365 993 399
rect 1061 365 1077 399
rect 1135 365 1151 399
rect 1219 365 1235 399
rect 1293 365 1309 399
rect 1377 365 1393 399
rect 1451 365 1467 399
rect 1535 365 1551 399
rect 1609 365 1625 399
rect 1693 365 1709 399
rect 1767 365 1783 399
rect 1851 365 1867 399
rect 1925 365 1941 399
rect 2009 365 2025 399
rect 2083 365 2099 399
rect 2167 365 2183 399
rect -2229 306 -2195 322
rect -2229 114 -2195 130
rect -2071 306 -2037 322
rect -2071 114 -2037 130
rect -1913 306 -1879 322
rect -1913 114 -1879 130
rect -1755 306 -1721 322
rect -1755 114 -1721 130
rect -1597 306 -1563 322
rect -1597 114 -1563 130
rect -1439 306 -1405 322
rect -1439 114 -1405 130
rect -1281 306 -1247 322
rect -1281 114 -1247 130
rect -1123 306 -1089 322
rect -1123 114 -1089 130
rect -965 306 -931 322
rect -965 114 -931 130
rect -807 306 -773 322
rect -807 114 -773 130
rect -649 306 -615 322
rect -649 114 -615 130
rect -491 306 -457 322
rect -491 114 -457 130
rect -333 306 -299 322
rect -333 114 -299 130
rect -175 306 -141 322
rect -175 114 -141 130
rect -17 306 17 322
rect -17 114 17 130
rect 141 306 175 322
rect 141 114 175 130
rect 299 306 333 322
rect 299 114 333 130
rect 457 306 491 322
rect 457 114 491 130
rect 615 306 649 322
rect 615 114 649 130
rect 773 306 807 322
rect 773 114 807 130
rect 931 306 965 322
rect 931 114 965 130
rect 1089 306 1123 322
rect 1089 114 1123 130
rect 1247 306 1281 322
rect 1247 114 1281 130
rect 1405 306 1439 322
rect 1405 114 1439 130
rect 1563 306 1597 322
rect 1563 114 1597 130
rect 1721 306 1755 322
rect 1721 114 1755 130
rect 1879 306 1913 322
rect 1879 114 1913 130
rect 2037 306 2071 322
rect 2037 114 2071 130
rect 2195 306 2229 322
rect 2195 114 2229 130
rect -2183 37 -2167 71
rect -2099 37 -2083 71
rect -2025 37 -2009 71
rect -1941 37 -1925 71
rect -1867 37 -1851 71
rect -1783 37 -1767 71
rect -1709 37 -1693 71
rect -1625 37 -1609 71
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -919 37 -903 71
rect -835 37 -819 71
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect 819 37 835 71
rect 903 37 919 71
rect 977 37 993 71
rect 1061 37 1077 71
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1609 37 1625 71
rect 1693 37 1709 71
rect 1767 37 1783 71
rect 1851 37 1867 71
rect 1925 37 1941 71
rect 2009 37 2025 71
rect 2083 37 2099 71
rect 2167 37 2183 71
rect -2183 -71 -2167 -37
rect -2099 -71 -2083 -37
rect -2025 -71 -2009 -37
rect -1941 -71 -1925 -37
rect -1867 -71 -1851 -37
rect -1783 -71 -1767 -37
rect -1709 -71 -1693 -37
rect -1625 -71 -1609 -37
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1609 -71 1625 -37
rect 1693 -71 1709 -37
rect 1767 -71 1783 -37
rect 1851 -71 1867 -37
rect 1925 -71 1941 -37
rect 2009 -71 2025 -37
rect 2083 -71 2099 -37
rect 2167 -71 2183 -37
rect -2229 -130 -2195 -114
rect -2229 -322 -2195 -306
rect -2071 -130 -2037 -114
rect -2071 -322 -2037 -306
rect -1913 -130 -1879 -114
rect -1913 -322 -1879 -306
rect -1755 -130 -1721 -114
rect -1755 -322 -1721 -306
rect -1597 -130 -1563 -114
rect -1597 -322 -1563 -306
rect -1439 -130 -1405 -114
rect -1439 -322 -1405 -306
rect -1281 -130 -1247 -114
rect -1281 -322 -1247 -306
rect -1123 -130 -1089 -114
rect -1123 -322 -1089 -306
rect -965 -130 -931 -114
rect -965 -322 -931 -306
rect -807 -130 -773 -114
rect -807 -322 -773 -306
rect -649 -130 -615 -114
rect -649 -322 -615 -306
rect -491 -130 -457 -114
rect -491 -322 -457 -306
rect -333 -130 -299 -114
rect -333 -322 -299 -306
rect -175 -130 -141 -114
rect -175 -322 -141 -306
rect -17 -130 17 -114
rect -17 -322 17 -306
rect 141 -130 175 -114
rect 141 -322 175 -306
rect 299 -130 333 -114
rect 299 -322 333 -306
rect 457 -130 491 -114
rect 457 -322 491 -306
rect 615 -130 649 -114
rect 615 -322 649 -306
rect 773 -130 807 -114
rect 773 -322 807 -306
rect 931 -130 965 -114
rect 931 -322 965 -306
rect 1089 -130 1123 -114
rect 1089 -322 1123 -306
rect 1247 -130 1281 -114
rect 1247 -322 1281 -306
rect 1405 -130 1439 -114
rect 1405 -322 1439 -306
rect 1563 -130 1597 -114
rect 1563 -322 1597 -306
rect 1721 -130 1755 -114
rect 1721 -322 1755 -306
rect 1879 -130 1913 -114
rect 1879 -322 1913 -306
rect 2037 -130 2071 -114
rect 2037 -322 2071 -306
rect 2195 -130 2229 -114
rect 2195 -322 2229 -306
rect -2183 -399 -2167 -365
rect -2099 -399 -2083 -365
rect -2025 -399 -2009 -365
rect -1941 -399 -1925 -365
rect -1867 -399 -1851 -365
rect -1783 -399 -1767 -365
rect -1709 -399 -1693 -365
rect -1625 -399 -1609 -365
rect -1551 -399 -1535 -365
rect -1467 -399 -1451 -365
rect -1393 -399 -1377 -365
rect -1309 -399 -1293 -365
rect -1235 -399 -1219 -365
rect -1151 -399 -1135 -365
rect -1077 -399 -1061 -365
rect -993 -399 -977 -365
rect -919 -399 -903 -365
rect -835 -399 -819 -365
rect -761 -399 -745 -365
rect -677 -399 -661 -365
rect -603 -399 -587 -365
rect -519 -399 -503 -365
rect -445 -399 -429 -365
rect -361 -399 -345 -365
rect -287 -399 -271 -365
rect -203 -399 -187 -365
rect -129 -399 -113 -365
rect -45 -399 -29 -365
rect 29 -399 45 -365
rect 113 -399 129 -365
rect 187 -399 203 -365
rect 271 -399 287 -365
rect 345 -399 361 -365
rect 429 -399 445 -365
rect 503 -399 519 -365
rect 587 -399 603 -365
rect 661 -399 677 -365
rect 745 -399 761 -365
rect 819 -399 835 -365
rect 903 -399 919 -365
rect 977 -399 993 -365
rect 1061 -399 1077 -365
rect 1135 -399 1151 -365
rect 1219 -399 1235 -365
rect 1293 -399 1309 -365
rect 1377 -399 1393 -365
rect 1451 -399 1467 -365
rect 1535 -399 1551 -365
rect 1609 -399 1625 -365
rect 1693 -399 1709 -365
rect 1767 -399 1783 -365
rect 1851 -399 1867 -365
rect 1925 -399 1941 -365
rect 2009 -399 2025 -365
rect 2083 -399 2099 -365
rect 2167 -399 2183 -365
rect -2183 -507 -2167 -473
rect -2099 -507 -2083 -473
rect -2025 -507 -2009 -473
rect -1941 -507 -1925 -473
rect -1867 -507 -1851 -473
rect -1783 -507 -1767 -473
rect -1709 -507 -1693 -473
rect -1625 -507 -1609 -473
rect -1551 -507 -1535 -473
rect -1467 -507 -1451 -473
rect -1393 -507 -1377 -473
rect -1309 -507 -1293 -473
rect -1235 -507 -1219 -473
rect -1151 -507 -1135 -473
rect -1077 -507 -1061 -473
rect -993 -507 -977 -473
rect -919 -507 -903 -473
rect -835 -507 -819 -473
rect -761 -507 -745 -473
rect -677 -507 -661 -473
rect -603 -507 -587 -473
rect -519 -507 -503 -473
rect -445 -507 -429 -473
rect -361 -507 -345 -473
rect -287 -507 -271 -473
rect -203 -507 -187 -473
rect -129 -507 -113 -473
rect -45 -507 -29 -473
rect 29 -507 45 -473
rect 113 -507 129 -473
rect 187 -507 203 -473
rect 271 -507 287 -473
rect 345 -507 361 -473
rect 429 -507 445 -473
rect 503 -507 519 -473
rect 587 -507 603 -473
rect 661 -507 677 -473
rect 745 -507 761 -473
rect 819 -507 835 -473
rect 903 -507 919 -473
rect 977 -507 993 -473
rect 1061 -507 1077 -473
rect 1135 -507 1151 -473
rect 1219 -507 1235 -473
rect 1293 -507 1309 -473
rect 1377 -507 1393 -473
rect 1451 -507 1467 -473
rect 1535 -507 1551 -473
rect 1609 -507 1625 -473
rect 1693 -507 1709 -473
rect 1767 -507 1783 -473
rect 1851 -507 1867 -473
rect 1925 -507 1941 -473
rect 2009 -507 2025 -473
rect 2083 -507 2099 -473
rect 2167 -507 2183 -473
rect -2229 -566 -2195 -550
rect -2229 -758 -2195 -742
rect -2071 -566 -2037 -550
rect -2071 -758 -2037 -742
rect -1913 -566 -1879 -550
rect -1913 -758 -1879 -742
rect -1755 -566 -1721 -550
rect -1755 -758 -1721 -742
rect -1597 -566 -1563 -550
rect -1597 -758 -1563 -742
rect -1439 -566 -1405 -550
rect -1439 -758 -1405 -742
rect -1281 -566 -1247 -550
rect -1281 -758 -1247 -742
rect -1123 -566 -1089 -550
rect -1123 -758 -1089 -742
rect -965 -566 -931 -550
rect -965 -758 -931 -742
rect -807 -566 -773 -550
rect -807 -758 -773 -742
rect -649 -566 -615 -550
rect -649 -758 -615 -742
rect -491 -566 -457 -550
rect -491 -758 -457 -742
rect -333 -566 -299 -550
rect -333 -758 -299 -742
rect -175 -566 -141 -550
rect -175 -758 -141 -742
rect -17 -566 17 -550
rect -17 -758 17 -742
rect 141 -566 175 -550
rect 141 -758 175 -742
rect 299 -566 333 -550
rect 299 -758 333 -742
rect 457 -566 491 -550
rect 457 -758 491 -742
rect 615 -566 649 -550
rect 615 -758 649 -742
rect 773 -566 807 -550
rect 773 -758 807 -742
rect 931 -566 965 -550
rect 931 -758 965 -742
rect 1089 -566 1123 -550
rect 1089 -758 1123 -742
rect 1247 -566 1281 -550
rect 1247 -758 1281 -742
rect 1405 -566 1439 -550
rect 1405 -758 1439 -742
rect 1563 -566 1597 -550
rect 1563 -758 1597 -742
rect 1721 -566 1755 -550
rect 1721 -758 1755 -742
rect 1879 -566 1913 -550
rect 1879 -758 1913 -742
rect 2037 -566 2071 -550
rect 2037 -758 2071 -742
rect 2195 -566 2229 -550
rect 2195 -758 2229 -742
rect -2183 -835 -2167 -801
rect -2099 -835 -2083 -801
rect -2025 -835 -2009 -801
rect -1941 -835 -1925 -801
rect -1867 -835 -1851 -801
rect -1783 -835 -1767 -801
rect -1709 -835 -1693 -801
rect -1625 -835 -1609 -801
rect -1551 -835 -1535 -801
rect -1467 -835 -1451 -801
rect -1393 -835 -1377 -801
rect -1309 -835 -1293 -801
rect -1235 -835 -1219 -801
rect -1151 -835 -1135 -801
rect -1077 -835 -1061 -801
rect -993 -835 -977 -801
rect -919 -835 -903 -801
rect -835 -835 -819 -801
rect -761 -835 -745 -801
rect -677 -835 -661 -801
rect -603 -835 -587 -801
rect -519 -835 -503 -801
rect -445 -835 -429 -801
rect -361 -835 -345 -801
rect -287 -835 -271 -801
rect -203 -835 -187 -801
rect -129 -835 -113 -801
rect -45 -835 -29 -801
rect 29 -835 45 -801
rect 113 -835 129 -801
rect 187 -835 203 -801
rect 271 -835 287 -801
rect 345 -835 361 -801
rect 429 -835 445 -801
rect 503 -835 519 -801
rect 587 -835 603 -801
rect 661 -835 677 -801
rect 745 -835 761 -801
rect 819 -835 835 -801
rect 903 -835 919 -801
rect 977 -835 993 -801
rect 1061 -835 1077 -801
rect 1135 -835 1151 -801
rect 1219 -835 1235 -801
rect 1293 -835 1309 -801
rect 1377 -835 1393 -801
rect 1451 -835 1467 -801
rect 1535 -835 1551 -801
rect 1609 -835 1625 -801
rect 1693 -835 1709 -801
rect 1767 -835 1783 -801
rect 1851 -835 1867 -801
rect 1925 -835 1941 -801
rect 2009 -835 2025 -801
rect 2083 -835 2099 -801
rect 2167 -835 2183 -801
rect -2183 -943 -2167 -909
rect -2099 -943 -2083 -909
rect -2025 -943 -2009 -909
rect -1941 -943 -1925 -909
rect -1867 -943 -1851 -909
rect -1783 -943 -1767 -909
rect -1709 -943 -1693 -909
rect -1625 -943 -1609 -909
rect -1551 -943 -1535 -909
rect -1467 -943 -1451 -909
rect -1393 -943 -1377 -909
rect -1309 -943 -1293 -909
rect -1235 -943 -1219 -909
rect -1151 -943 -1135 -909
rect -1077 -943 -1061 -909
rect -993 -943 -977 -909
rect -919 -943 -903 -909
rect -835 -943 -819 -909
rect -761 -943 -745 -909
rect -677 -943 -661 -909
rect -603 -943 -587 -909
rect -519 -943 -503 -909
rect -445 -943 -429 -909
rect -361 -943 -345 -909
rect -287 -943 -271 -909
rect -203 -943 -187 -909
rect -129 -943 -113 -909
rect -45 -943 -29 -909
rect 29 -943 45 -909
rect 113 -943 129 -909
rect 187 -943 203 -909
rect 271 -943 287 -909
rect 345 -943 361 -909
rect 429 -943 445 -909
rect 503 -943 519 -909
rect 587 -943 603 -909
rect 661 -943 677 -909
rect 745 -943 761 -909
rect 819 -943 835 -909
rect 903 -943 919 -909
rect 977 -943 993 -909
rect 1061 -943 1077 -909
rect 1135 -943 1151 -909
rect 1219 -943 1235 -909
rect 1293 -943 1309 -909
rect 1377 -943 1393 -909
rect 1451 -943 1467 -909
rect 1535 -943 1551 -909
rect 1609 -943 1625 -909
rect 1693 -943 1709 -909
rect 1767 -943 1783 -909
rect 1851 -943 1867 -909
rect 1925 -943 1941 -909
rect 2009 -943 2025 -909
rect 2083 -943 2099 -909
rect 2167 -943 2183 -909
rect -2229 -1002 -2195 -986
rect -2229 -1194 -2195 -1178
rect -2071 -1002 -2037 -986
rect -2071 -1194 -2037 -1178
rect -1913 -1002 -1879 -986
rect -1913 -1194 -1879 -1178
rect -1755 -1002 -1721 -986
rect -1755 -1194 -1721 -1178
rect -1597 -1002 -1563 -986
rect -1597 -1194 -1563 -1178
rect -1439 -1002 -1405 -986
rect -1439 -1194 -1405 -1178
rect -1281 -1002 -1247 -986
rect -1281 -1194 -1247 -1178
rect -1123 -1002 -1089 -986
rect -1123 -1194 -1089 -1178
rect -965 -1002 -931 -986
rect -965 -1194 -931 -1178
rect -807 -1002 -773 -986
rect -807 -1194 -773 -1178
rect -649 -1002 -615 -986
rect -649 -1194 -615 -1178
rect -491 -1002 -457 -986
rect -491 -1194 -457 -1178
rect -333 -1002 -299 -986
rect -333 -1194 -299 -1178
rect -175 -1002 -141 -986
rect -175 -1194 -141 -1178
rect -17 -1002 17 -986
rect -17 -1194 17 -1178
rect 141 -1002 175 -986
rect 141 -1194 175 -1178
rect 299 -1002 333 -986
rect 299 -1194 333 -1178
rect 457 -1002 491 -986
rect 457 -1194 491 -1178
rect 615 -1002 649 -986
rect 615 -1194 649 -1178
rect 773 -1002 807 -986
rect 773 -1194 807 -1178
rect 931 -1002 965 -986
rect 931 -1194 965 -1178
rect 1089 -1002 1123 -986
rect 1089 -1194 1123 -1178
rect 1247 -1002 1281 -986
rect 1247 -1194 1281 -1178
rect 1405 -1002 1439 -986
rect 1405 -1194 1439 -1178
rect 1563 -1002 1597 -986
rect 1563 -1194 1597 -1178
rect 1721 -1002 1755 -986
rect 1721 -1194 1755 -1178
rect 1879 -1002 1913 -986
rect 1879 -1194 1913 -1178
rect 2037 -1002 2071 -986
rect 2037 -1194 2071 -1178
rect 2195 -1002 2229 -986
rect 2195 -1194 2229 -1178
rect -2183 -1271 -2167 -1237
rect -2099 -1271 -2083 -1237
rect -2025 -1271 -2009 -1237
rect -1941 -1271 -1925 -1237
rect -1867 -1271 -1851 -1237
rect -1783 -1271 -1767 -1237
rect -1709 -1271 -1693 -1237
rect -1625 -1271 -1609 -1237
rect -1551 -1271 -1535 -1237
rect -1467 -1271 -1451 -1237
rect -1393 -1271 -1377 -1237
rect -1309 -1271 -1293 -1237
rect -1235 -1271 -1219 -1237
rect -1151 -1271 -1135 -1237
rect -1077 -1271 -1061 -1237
rect -993 -1271 -977 -1237
rect -919 -1271 -903 -1237
rect -835 -1271 -819 -1237
rect -761 -1271 -745 -1237
rect -677 -1271 -661 -1237
rect -603 -1271 -587 -1237
rect -519 -1271 -503 -1237
rect -445 -1271 -429 -1237
rect -361 -1271 -345 -1237
rect -287 -1271 -271 -1237
rect -203 -1271 -187 -1237
rect -129 -1271 -113 -1237
rect -45 -1271 -29 -1237
rect 29 -1271 45 -1237
rect 113 -1271 129 -1237
rect 187 -1271 203 -1237
rect 271 -1271 287 -1237
rect 345 -1271 361 -1237
rect 429 -1271 445 -1237
rect 503 -1271 519 -1237
rect 587 -1271 603 -1237
rect 661 -1271 677 -1237
rect 745 -1271 761 -1237
rect 819 -1271 835 -1237
rect 903 -1271 919 -1237
rect 977 -1271 993 -1237
rect 1061 -1271 1077 -1237
rect 1135 -1271 1151 -1237
rect 1219 -1271 1235 -1237
rect 1293 -1271 1309 -1237
rect 1377 -1271 1393 -1237
rect 1451 -1271 1467 -1237
rect 1535 -1271 1551 -1237
rect 1609 -1271 1625 -1237
rect 1693 -1271 1709 -1237
rect 1767 -1271 1783 -1237
rect 1851 -1271 1867 -1237
rect 1925 -1271 1941 -1237
rect 2009 -1271 2025 -1237
rect 2083 -1271 2099 -1237
rect 2167 -1271 2183 -1237
rect -2183 -1379 -2167 -1345
rect -2099 -1379 -2083 -1345
rect -2025 -1379 -2009 -1345
rect -1941 -1379 -1925 -1345
rect -1867 -1379 -1851 -1345
rect -1783 -1379 -1767 -1345
rect -1709 -1379 -1693 -1345
rect -1625 -1379 -1609 -1345
rect -1551 -1379 -1535 -1345
rect -1467 -1379 -1451 -1345
rect -1393 -1379 -1377 -1345
rect -1309 -1379 -1293 -1345
rect -1235 -1379 -1219 -1345
rect -1151 -1379 -1135 -1345
rect -1077 -1379 -1061 -1345
rect -993 -1379 -977 -1345
rect -919 -1379 -903 -1345
rect -835 -1379 -819 -1345
rect -761 -1379 -745 -1345
rect -677 -1379 -661 -1345
rect -603 -1379 -587 -1345
rect -519 -1379 -503 -1345
rect -445 -1379 -429 -1345
rect -361 -1379 -345 -1345
rect -287 -1379 -271 -1345
rect -203 -1379 -187 -1345
rect -129 -1379 -113 -1345
rect -45 -1379 -29 -1345
rect 29 -1379 45 -1345
rect 113 -1379 129 -1345
rect 187 -1379 203 -1345
rect 271 -1379 287 -1345
rect 345 -1379 361 -1345
rect 429 -1379 445 -1345
rect 503 -1379 519 -1345
rect 587 -1379 603 -1345
rect 661 -1379 677 -1345
rect 745 -1379 761 -1345
rect 819 -1379 835 -1345
rect 903 -1379 919 -1345
rect 977 -1379 993 -1345
rect 1061 -1379 1077 -1345
rect 1135 -1379 1151 -1345
rect 1219 -1379 1235 -1345
rect 1293 -1379 1309 -1345
rect 1377 -1379 1393 -1345
rect 1451 -1379 1467 -1345
rect 1535 -1379 1551 -1345
rect 1609 -1379 1625 -1345
rect 1693 -1379 1709 -1345
rect 1767 -1379 1783 -1345
rect 1851 -1379 1867 -1345
rect 1925 -1379 1941 -1345
rect 2009 -1379 2025 -1345
rect 2083 -1379 2099 -1345
rect 2167 -1379 2183 -1345
rect -2229 -1438 -2195 -1422
rect -2229 -1630 -2195 -1614
rect -2071 -1438 -2037 -1422
rect -2071 -1630 -2037 -1614
rect -1913 -1438 -1879 -1422
rect -1913 -1630 -1879 -1614
rect -1755 -1438 -1721 -1422
rect -1755 -1630 -1721 -1614
rect -1597 -1438 -1563 -1422
rect -1597 -1630 -1563 -1614
rect -1439 -1438 -1405 -1422
rect -1439 -1630 -1405 -1614
rect -1281 -1438 -1247 -1422
rect -1281 -1630 -1247 -1614
rect -1123 -1438 -1089 -1422
rect -1123 -1630 -1089 -1614
rect -965 -1438 -931 -1422
rect -965 -1630 -931 -1614
rect -807 -1438 -773 -1422
rect -807 -1630 -773 -1614
rect -649 -1438 -615 -1422
rect -649 -1630 -615 -1614
rect -491 -1438 -457 -1422
rect -491 -1630 -457 -1614
rect -333 -1438 -299 -1422
rect -333 -1630 -299 -1614
rect -175 -1438 -141 -1422
rect -175 -1630 -141 -1614
rect -17 -1438 17 -1422
rect -17 -1630 17 -1614
rect 141 -1438 175 -1422
rect 141 -1630 175 -1614
rect 299 -1438 333 -1422
rect 299 -1630 333 -1614
rect 457 -1438 491 -1422
rect 457 -1630 491 -1614
rect 615 -1438 649 -1422
rect 615 -1630 649 -1614
rect 773 -1438 807 -1422
rect 773 -1630 807 -1614
rect 931 -1438 965 -1422
rect 931 -1630 965 -1614
rect 1089 -1438 1123 -1422
rect 1089 -1630 1123 -1614
rect 1247 -1438 1281 -1422
rect 1247 -1630 1281 -1614
rect 1405 -1438 1439 -1422
rect 1405 -1630 1439 -1614
rect 1563 -1438 1597 -1422
rect 1563 -1630 1597 -1614
rect 1721 -1438 1755 -1422
rect 1721 -1630 1755 -1614
rect 1879 -1438 1913 -1422
rect 1879 -1630 1913 -1614
rect 2037 -1438 2071 -1422
rect 2037 -1630 2071 -1614
rect 2195 -1438 2229 -1422
rect 2195 -1630 2229 -1614
rect -2183 -1707 -2167 -1673
rect -2099 -1707 -2083 -1673
rect -2025 -1707 -2009 -1673
rect -1941 -1707 -1925 -1673
rect -1867 -1707 -1851 -1673
rect -1783 -1707 -1767 -1673
rect -1709 -1707 -1693 -1673
rect -1625 -1707 -1609 -1673
rect -1551 -1707 -1535 -1673
rect -1467 -1707 -1451 -1673
rect -1393 -1707 -1377 -1673
rect -1309 -1707 -1293 -1673
rect -1235 -1707 -1219 -1673
rect -1151 -1707 -1135 -1673
rect -1077 -1707 -1061 -1673
rect -993 -1707 -977 -1673
rect -919 -1707 -903 -1673
rect -835 -1707 -819 -1673
rect -761 -1707 -745 -1673
rect -677 -1707 -661 -1673
rect -603 -1707 -587 -1673
rect -519 -1707 -503 -1673
rect -445 -1707 -429 -1673
rect -361 -1707 -345 -1673
rect -287 -1707 -271 -1673
rect -203 -1707 -187 -1673
rect -129 -1707 -113 -1673
rect -45 -1707 -29 -1673
rect 29 -1707 45 -1673
rect 113 -1707 129 -1673
rect 187 -1707 203 -1673
rect 271 -1707 287 -1673
rect 345 -1707 361 -1673
rect 429 -1707 445 -1673
rect 503 -1707 519 -1673
rect 587 -1707 603 -1673
rect 661 -1707 677 -1673
rect 745 -1707 761 -1673
rect 819 -1707 835 -1673
rect 903 -1707 919 -1673
rect 977 -1707 993 -1673
rect 1061 -1707 1077 -1673
rect 1135 -1707 1151 -1673
rect 1219 -1707 1235 -1673
rect 1293 -1707 1309 -1673
rect 1377 -1707 1393 -1673
rect 1451 -1707 1467 -1673
rect 1535 -1707 1551 -1673
rect 1609 -1707 1625 -1673
rect 1693 -1707 1709 -1673
rect 1767 -1707 1783 -1673
rect 1851 -1707 1867 -1673
rect 1925 -1707 1941 -1673
rect 2009 -1707 2025 -1673
rect 2083 -1707 2099 -1673
rect 2167 -1707 2183 -1673
rect -2183 -1815 -2167 -1781
rect -2099 -1815 -2083 -1781
rect -2025 -1815 -2009 -1781
rect -1941 -1815 -1925 -1781
rect -1867 -1815 -1851 -1781
rect -1783 -1815 -1767 -1781
rect -1709 -1815 -1693 -1781
rect -1625 -1815 -1609 -1781
rect -1551 -1815 -1535 -1781
rect -1467 -1815 -1451 -1781
rect -1393 -1815 -1377 -1781
rect -1309 -1815 -1293 -1781
rect -1235 -1815 -1219 -1781
rect -1151 -1815 -1135 -1781
rect -1077 -1815 -1061 -1781
rect -993 -1815 -977 -1781
rect -919 -1815 -903 -1781
rect -835 -1815 -819 -1781
rect -761 -1815 -745 -1781
rect -677 -1815 -661 -1781
rect -603 -1815 -587 -1781
rect -519 -1815 -503 -1781
rect -445 -1815 -429 -1781
rect -361 -1815 -345 -1781
rect -287 -1815 -271 -1781
rect -203 -1815 -187 -1781
rect -129 -1815 -113 -1781
rect -45 -1815 -29 -1781
rect 29 -1815 45 -1781
rect 113 -1815 129 -1781
rect 187 -1815 203 -1781
rect 271 -1815 287 -1781
rect 345 -1815 361 -1781
rect 429 -1815 445 -1781
rect 503 -1815 519 -1781
rect 587 -1815 603 -1781
rect 661 -1815 677 -1781
rect 745 -1815 761 -1781
rect 819 -1815 835 -1781
rect 903 -1815 919 -1781
rect 977 -1815 993 -1781
rect 1061 -1815 1077 -1781
rect 1135 -1815 1151 -1781
rect 1219 -1815 1235 -1781
rect 1293 -1815 1309 -1781
rect 1377 -1815 1393 -1781
rect 1451 -1815 1467 -1781
rect 1535 -1815 1551 -1781
rect 1609 -1815 1625 -1781
rect 1693 -1815 1709 -1781
rect 1767 -1815 1783 -1781
rect 1851 -1815 1867 -1781
rect 1925 -1815 1941 -1781
rect 2009 -1815 2025 -1781
rect 2083 -1815 2099 -1781
rect 2167 -1815 2183 -1781
rect -2229 -1874 -2195 -1858
rect -2229 -2066 -2195 -2050
rect -2071 -1874 -2037 -1858
rect -2071 -2066 -2037 -2050
rect -1913 -1874 -1879 -1858
rect -1913 -2066 -1879 -2050
rect -1755 -1874 -1721 -1858
rect -1755 -2066 -1721 -2050
rect -1597 -1874 -1563 -1858
rect -1597 -2066 -1563 -2050
rect -1439 -1874 -1405 -1858
rect -1439 -2066 -1405 -2050
rect -1281 -1874 -1247 -1858
rect -1281 -2066 -1247 -2050
rect -1123 -1874 -1089 -1858
rect -1123 -2066 -1089 -2050
rect -965 -1874 -931 -1858
rect -965 -2066 -931 -2050
rect -807 -1874 -773 -1858
rect -807 -2066 -773 -2050
rect -649 -1874 -615 -1858
rect -649 -2066 -615 -2050
rect -491 -1874 -457 -1858
rect -491 -2066 -457 -2050
rect -333 -1874 -299 -1858
rect -333 -2066 -299 -2050
rect -175 -1874 -141 -1858
rect -175 -2066 -141 -2050
rect -17 -1874 17 -1858
rect -17 -2066 17 -2050
rect 141 -1874 175 -1858
rect 141 -2066 175 -2050
rect 299 -1874 333 -1858
rect 299 -2066 333 -2050
rect 457 -1874 491 -1858
rect 457 -2066 491 -2050
rect 615 -1874 649 -1858
rect 615 -2066 649 -2050
rect 773 -1874 807 -1858
rect 773 -2066 807 -2050
rect 931 -1874 965 -1858
rect 931 -2066 965 -2050
rect 1089 -1874 1123 -1858
rect 1089 -2066 1123 -2050
rect 1247 -1874 1281 -1858
rect 1247 -2066 1281 -2050
rect 1405 -1874 1439 -1858
rect 1405 -2066 1439 -2050
rect 1563 -1874 1597 -1858
rect 1563 -2066 1597 -2050
rect 1721 -1874 1755 -1858
rect 1721 -2066 1755 -2050
rect 1879 -1874 1913 -1858
rect 1879 -2066 1913 -2050
rect 2037 -1874 2071 -1858
rect 2037 -2066 2071 -2050
rect 2195 -1874 2229 -1858
rect 2195 -2066 2229 -2050
rect -2183 -2143 -2167 -2109
rect -2099 -2143 -2083 -2109
rect -2025 -2143 -2009 -2109
rect -1941 -2143 -1925 -2109
rect -1867 -2143 -1851 -2109
rect -1783 -2143 -1767 -2109
rect -1709 -2143 -1693 -2109
rect -1625 -2143 -1609 -2109
rect -1551 -2143 -1535 -2109
rect -1467 -2143 -1451 -2109
rect -1393 -2143 -1377 -2109
rect -1309 -2143 -1293 -2109
rect -1235 -2143 -1219 -2109
rect -1151 -2143 -1135 -2109
rect -1077 -2143 -1061 -2109
rect -993 -2143 -977 -2109
rect -919 -2143 -903 -2109
rect -835 -2143 -819 -2109
rect -761 -2143 -745 -2109
rect -677 -2143 -661 -2109
rect -603 -2143 -587 -2109
rect -519 -2143 -503 -2109
rect -445 -2143 -429 -2109
rect -361 -2143 -345 -2109
rect -287 -2143 -271 -2109
rect -203 -2143 -187 -2109
rect -129 -2143 -113 -2109
rect -45 -2143 -29 -2109
rect 29 -2143 45 -2109
rect 113 -2143 129 -2109
rect 187 -2143 203 -2109
rect 271 -2143 287 -2109
rect 345 -2143 361 -2109
rect 429 -2143 445 -2109
rect 503 -2143 519 -2109
rect 587 -2143 603 -2109
rect 661 -2143 677 -2109
rect 745 -2143 761 -2109
rect 819 -2143 835 -2109
rect 903 -2143 919 -2109
rect 977 -2143 993 -2109
rect 1061 -2143 1077 -2109
rect 1135 -2143 1151 -2109
rect 1219 -2143 1235 -2109
rect 1293 -2143 1309 -2109
rect 1377 -2143 1393 -2109
rect 1451 -2143 1467 -2109
rect 1535 -2143 1551 -2109
rect 1609 -2143 1625 -2109
rect 1693 -2143 1709 -2109
rect 1767 -2143 1783 -2109
rect 1851 -2143 1867 -2109
rect 1925 -2143 1941 -2109
rect 2009 -2143 2025 -2109
rect 2083 -2143 2099 -2109
rect 2167 -2143 2183 -2109
rect -2363 -2247 -2329 -2185
rect 2329 -2247 2363 -2185
rect -2363 -2281 -2267 -2247
rect 2267 -2281 2363 -2247
<< viali >>
rect -2167 2109 -2099 2143
rect -2009 2109 -1941 2143
rect -1851 2109 -1783 2143
rect -1693 2109 -1625 2143
rect -1535 2109 -1467 2143
rect -1377 2109 -1309 2143
rect -1219 2109 -1151 2143
rect -1061 2109 -993 2143
rect -903 2109 -835 2143
rect -745 2109 -677 2143
rect -587 2109 -519 2143
rect -429 2109 -361 2143
rect -271 2109 -203 2143
rect -113 2109 -45 2143
rect 45 2109 113 2143
rect 203 2109 271 2143
rect 361 2109 429 2143
rect 519 2109 587 2143
rect 677 2109 745 2143
rect 835 2109 903 2143
rect 993 2109 1061 2143
rect 1151 2109 1219 2143
rect 1309 2109 1377 2143
rect 1467 2109 1535 2143
rect 1625 2109 1693 2143
rect 1783 2109 1851 2143
rect 1941 2109 2009 2143
rect 2099 2109 2167 2143
rect -2229 1874 -2195 2050
rect -2071 1874 -2037 2050
rect -1913 1874 -1879 2050
rect -1755 1874 -1721 2050
rect -1597 1874 -1563 2050
rect -1439 1874 -1405 2050
rect -1281 1874 -1247 2050
rect -1123 1874 -1089 2050
rect -965 1874 -931 2050
rect -807 1874 -773 2050
rect -649 1874 -615 2050
rect -491 1874 -457 2050
rect -333 1874 -299 2050
rect -175 1874 -141 2050
rect -17 1874 17 2050
rect 141 1874 175 2050
rect 299 1874 333 2050
rect 457 1874 491 2050
rect 615 1874 649 2050
rect 773 1874 807 2050
rect 931 1874 965 2050
rect 1089 1874 1123 2050
rect 1247 1874 1281 2050
rect 1405 1874 1439 2050
rect 1563 1874 1597 2050
rect 1721 1874 1755 2050
rect 1879 1874 1913 2050
rect 2037 1874 2071 2050
rect 2195 1874 2229 2050
rect -2167 1781 -2099 1815
rect -2009 1781 -1941 1815
rect -1851 1781 -1783 1815
rect -1693 1781 -1625 1815
rect -1535 1781 -1467 1815
rect -1377 1781 -1309 1815
rect -1219 1781 -1151 1815
rect -1061 1781 -993 1815
rect -903 1781 -835 1815
rect -745 1781 -677 1815
rect -587 1781 -519 1815
rect -429 1781 -361 1815
rect -271 1781 -203 1815
rect -113 1781 -45 1815
rect 45 1781 113 1815
rect 203 1781 271 1815
rect 361 1781 429 1815
rect 519 1781 587 1815
rect 677 1781 745 1815
rect 835 1781 903 1815
rect 993 1781 1061 1815
rect 1151 1781 1219 1815
rect 1309 1781 1377 1815
rect 1467 1781 1535 1815
rect 1625 1781 1693 1815
rect 1783 1781 1851 1815
rect 1941 1781 2009 1815
rect 2099 1781 2167 1815
rect -2167 1673 -2099 1707
rect -2009 1673 -1941 1707
rect -1851 1673 -1783 1707
rect -1693 1673 -1625 1707
rect -1535 1673 -1467 1707
rect -1377 1673 -1309 1707
rect -1219 1673 -1151 1707
rect -1061 1673 -993 1707
rect -903 1673 -835 1707
rect -745 1673 -677 1707
rect -587 1673 -519 1707
rect -429 1673 -361 1707
rect -271 1673 -203 1707
rect -113 1673 -45 1707
rect 45 1673 113 1707
rect 203 1673 271 1707
rect 361 1673 429 1707
rect 519 1673 587 1707
rect 677 1673 745 1707
rect 835 1673 903 1707
rect 993 1673 1061 1707
rect 1151 1673 1219 1707
rect 1309 1673 1377 1707
rect 1467 1673 1535 1707
rect 1625 1673 1693 1707
rect 1783 1673 1851 1707
rect 1941 1673 2009 1707
rect 2099 1673 2167 1707
rect -2229 1438 -2195 1614
rect -2071 1438 -2037 1614
rect -1913 1438 -1879 1614
rect -1755 1438 -1721 1614
rect -1597 1438 -1563 1614
rect -1439 1438 -1405 1614
rect -1281 1438 -1247 1614
rect -1123 1438 -1089 1614
rect -965 1438 -931 1614
rect -807 1438 -773 1614
rect -649 1438 -615 1614
rect -491 1438 -457 1614
rect -333 1438 -299 1614
rect -175 1438 -141 1614
rect -17 1438 17 1614
rect 141 1438 175 1614
rect 299 1438 333 1614
rect 457 1438 491 1614
rect 615 1438 649 1614
rect 773 1438 807 1614
rect 931 1438 965 1614
rect 1089 1438 1123 1614
rect 1247 1438 1281 1614
rect 1405 1438 1439 1614
rect 1563 1438 1597 1614
rect 1721 1438 1755 1614
rect 1879 1438 1913 1614
rect 2037 1438 2071 1614
rect 2195 1438 2229 1614
rect -2167 1345 -2099 1379
rect -2009 1345 -1941 1379
rect -1851 1345 -1783 1379
rect -1693 1345 -1625 1379
rect -1535 1345 -1467 1379
rect -1377 1345 -1309 1379
rect -1219 1345 -1151 1379
rect -1061 1345 -993 1379
rect -903 1345 -835 1379
rect -745 1345 -677 1379
rect -587 1345 -519 1379
rect -429 1345 -361 1379
rect -271 1345 -203 1379
rect -113 1345 -45 1379
rect 45 1345 113 1379
rect 203 1345 271 1379
rect 361 1345 429 1379
rect 519 1345 587 1379
rect 677 1345 745 1379
rect 835 1345 903 1379
rect 993 1345 1061 1379
rect 1151 1345 1219 1379
rect 1309 1345 1377 1379
rect 1467 1345 1535 1379
rect 1625 1345 1693 1379
rect 1783 1345 1851 1379
rect 1941 1345 2009 1379
rect 2099 1345 2167 1379
rect -2167 1237 -2099 1271
rect -2009 1237 -1941 1271
rect -1851 1237 -1783 1271
rect -1693 1237 -1625 1271
rect -1535 1237 -1467 1271
rect -1377 1237 -1309 1271
rect -1219 1237 -1151 1271
rect -1061 1237 -993 1271
rect -903 1237 -835 1271
rect -745 1237 -677 1271
rect -587 1237 -519 1271
rect -429 1237 -361 1271
rect -271 1237 -203 1271
rect -113 1237 -45 1271
rect 45 1237 113 1271
rect 203 1237 271 1271
rect 361 1237 429 1271
rect 519 1237 587 1271
rect 677 1237 745 1271
rect 835 1237 903 1271
rect 993 1237 1061 1271
rect 1151 1237 1219 1271
rect 1309 1237 1377 1271
rect 1467 1237 1535 1271
rect 1625 1237 1693 1271
rect 1783 1237 1851 1271
rect 1941 1237 2009 1271
rect 2099 1237 2167 1271
rect -2229 1002 -2195 1178
rect -2071 1002 -2037 1178
rect -1913 1002 -1879 1178
rect -1755 1002 -1721 1178
rect -1597 1002 -1563 1178
rect -1439 1002 -1405 1178
rect -1281 1002 -1247 1178
rect -1123 1002 -1089 1178
rect -965 1002 -931 1178
rect -807 1002 -773 1178
rect -649 1002 -615 1178
rect -491 1002 -457 1178
rect -333 1002 -299 1178
rect -175 1002 -141 1178
rect -17 1002 17 1178
rect 141 1002 175 1178
rect 299 1002 333 1178
rect 457 1002 491 1178
rect 615 1002 649 1178
rect 773 1002 807 1178
rect 931 1002 965 1178
rect 1089 1002 1123 1178
rect 1247 1002 1281 1178
rect 1405 1002 1439 1178
rect 1563 1002 1597 1178
rect 1721 1002 1755 1178
rect 1879 1002 1913 1178
rect 2037 1002 2071 1178
rect 2195 1002 2229 1178
rect -2167 909 -2099 943
rect -2009 909 -1941 943
rect -1851 909 -1783 943
rect -1693 909 -1625 943
rect -1535 909 -1467 943
rect -1377 909 -1309 943
rect -1219 909 -1151 943
rect -1061 909 -993 943
rect -903 909 -835 943
rect -745 909 -677 943
rect -587 909 -519 943
rect -429 909 -361 943
rect -271 909 -203 943
rect -113 909 -45 943
rect 45 909 113 943
rect 203 909 271 943
rect 361 909 429 943
rect 519 909 587 943
rect 677 909 745 943
rect 835 909 903 943
rect 993 909 1061 943
rect 1151 909 1219 943
rect 1309 909 1377 943
rect 1467 909 1535 943
rect 1625 909 1693 943
rect 1783 909 1851 943
rect 1941 909 2009 943
rect 2099 909 2167 943
rect -2167 801 -2099 835
rect -2009 801 -1941 835
rect -1851 801 -1783 835
rect -1693 801 -1625 835
rect -1535 801 -1467 835
rect -1377 801 -1309 835
rect -1219 801 -1151 835
rect -1061 801 -993 835
rect -903 801 -835 835
rect -745 801 -677 835
rect -587 801 -519 835
rect -429 801 -361 835
rect -271 801 -203 835
rect -113 801 -45 835
rect 45 801 113 835
rect 203 801 271 835
rect 361 801 429 835
rect 519 801 587 835
rect 677 801 745 835
rect 835 801 903 835
rect 993 801 1061 835
rect 1151 801 1219 835
rect 1309 801 1377 835
rect 1467 801 1535 835
rect 1625 801 1693 835
rect 1783 801 1851 835
rect 1941 801 2009 835
rect 2099 801 2167 835
rect -2229 566 -2195 742
rect -2071 566 -2037 742
rect -1913 566 -1879 742
rect -1755 566 -1721 742
rect -1597 566 -1563 742
rect -1439 566 -1405 742
rect -1281 566 -1247 742
rect -1123 566 -1089 742
rect -965 566 -931 742
rect -807 566 -773 742
rect -649 566 -615 742
rect -491 566 -457 742
rect -333 566 -299 742
rect -175 566 -141 742
rect -17 566 17 742
rect 141 566 175 742
rect 299 566 333 742
rect 457 566 491 742
rect 615 566 649 742
rect 773 566 807 742
rect 931 566 965 742
rect 1089 566 1123 742
rect 1247 566 1281 742
rect 1405 566 1439 742
rect 1563 566 1597 742
rect 1721 566 1755 742
rect 1879 566 1913 742
rect 2037 566 2071 742
rect 2195 566 2229 742
rect -2167 473 -2099 507
rect -2009 473 -1941 507
rect -1851 473 -1783 507
rect -1693 473 -1625 507
rect -1535 473 -1467 507
rect -1377 473 -1309 507
rect -1219 473 -1151 507
rect -1061 473 -993 507
rect -903 473 -835 507
rect -745 473 -677 507
rect -587 473 -519 507
rect -429 473 -361 507
rect -271 473 -203 507
rect -113 473 -45 507
rect 45 473 113 507
rect 203 473 271 507
rect 361 473 429 507
rect 519 473 587 507
rect 677 473 745 507
rect 835 473 903 507
rect 993 473 1061 507
rect 1151 473 1219 507
rect 1309 473 1377 507
rect 1467 473 1535 507
rect 1625 473 1693 507
rect 1783 473 1851 507
rect 1941 473 2009 507
rect 2099 473 2167 507
rect -2167 365 -2099 399
rect -2009 365 -1941 399
rect -1851 365 -1783 399
rect -1693 365 -1625 399
rect -1535 365 -1467 399
rect -1377 365 -1309 399
rect -1219 365 -1151 399
rect -1061 365 -993 399
rect -903 365 -835 399
rect -745 365 -677 399
rect -587 365 -519 399
rect -429 365 -361 399
rect -271 365 -203 399
rect -113 365 -45 399
rect 45 365 113 399
rect 203 365 271 399
rect 361 365 429 399
rect 519 365 587 399
rect 677 365 745 399
rect 835 365 903 399
rect 993 365 1061 399
rect 1151 365 1219 399
rect 1309 365 1377 399
rect 1467 365 1535 399
rect 1625 365 1693 399
rect 1783 365 1851 399
rect 1941 365 2009 399
rect 2099 365 2167 399
rect -2229 130 -2195 306
rect -2071 130 -2037 306
rect -1913 130 -1879 306
rect -1755 130 -1721 306
rect -1597 130 -1563 306
rect -1439 130 -1405 306
rect -1281 130 -1247 306
rect -1123 130 -1089 306
rect -965 130 -931 306
rect -807 130 -773 306
rect -649 130 -615 306
rect -491 130 -457 306
rect -333 130 -299 306
rect -175 130 -141 306
rect -17 130 17 306
rect 141 130 175 306
rect 299 130 333 306
rect 457 130 491 306
rect 615 130 649 306
rect 773 130 807 306
rect 931 130 965 306
rect 1089 130 1123 306
rect 1247 130 1281 306
rect 1405 130 1439 306
rect 1563 130 1597 306
rect 1721 130 1755 306
rect 1879 130 1913 306
rect 2037 130 2071 306
rect 2195 130 2229 306
rect -2167 37 -2099 71
rect -2009 37 -1941 71
rect -1851 37 -1783 71
rect -1693 37 -1625 71
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect 1625 37 1693 71
rect 1783 37 1851 71
rect 1941 37 2009 71
rect 2099 37 2167 71
rect -2167 -71 -2099 -37
rect -2009 -71 -1941 -37
rect -1851 -71 -1783 -37
rect -1693 -71 -1625 -37
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect 1625 -71 1693 -37
rect 1783 -71 1851 -37
rect 1941 -71 2009 -37
rect 2099 -71 2167 -37
rect -2229 -306 -2195 -130
rect -2071 -306 -2037 -130
rect -1913 -306 -1879 -130
rect -1755 -306 -1721 -130
rect -1597 -306 -1563 -130
rect -1439 -306 -1405 -130
rect -1281 -306 -1247 -130
rect -1123 -306 -1089 -130
rect -965 -306 -931 -130
rect -807 -306 -773 -130
rect -649 -306 -615 -130
rect -491 -306 -457 -130
rect -333 -306 -299 -130
rect -175 -306 -141 -130
rect -17 -306 17 -130
rect 141 -306 175 -130
rect 299 -306 333 -130
rect 457 -306 491 -130
rect 615 -306 649 -130
rect 773 -306 807 -130
rect 931 -306 965 -130
rect 1089 -306 1123 -130
rect 1247 -306 1281 -130
rect 1405 -306 1439 -130
rect 1563 -306 1597 -130
rect 1721 -306 1755 -130
rect 1879 -306 1913 -130
rect 2037 -306 2071 -130
rect 2195 -306 2229 -130
rect -2167 -399 -2099 -365
rect -2009 -399 -1941 -365
rect -1851 -399 -1783 -365
rect -1693 -399 -1625 -365
rect -1535 -399 -1467 -365
rect -1377 -399 -1309 -365
rect -1219 -399 -1151 -365
rect -1061 -399 -993 -365
rect -903 -399 -835 -365
rect -745 -399 -677 -365
rect -587 -399 -519 -365
rect -429 -399 -361 -365
rect -271 -399 -203 -365
rect -113 -399 -45 -365
rect 45 -399 113 -365
rect 203 -399 271 -365
rect 361 -399 429 -365
rect 519 -399 587 -365
rect 677 -399 745 -365
rect 835 -399 903 -365
rect 993 -399 1061 -365
rect 1151 -399 1219 -365
rect 1309 -399 1377 -365
rect 1467 -399 1535 -365
rect 1625 -399 1693 -365
rect 1783 -399 1851 -365
rect 1941 -399 2009 -365
rect 2099 -399 2167 -365
rect -2167 -507 -2099 -473
rect -2009 -507 -1941 -473
rect -1851 -507 -1783 -473
rect -1693 -507 -1625 -473
rect -1535 -507 -1467 -473
rect -1377 -507 -1309 -473
rect -1219 -507 -1151 -473
rect -1061 -507 -993 -473
rect -903 -507 -835 -473
rect -745 -507 -677 -473
rect -587 -507 -519 -473
rect -429 -507 -361 -473
rect -271 -507 -203 -473
rect -113 -507 -45 -473
rect 45 -507 113 -473
rect 203 -507 271 -473
rect 361 -507 429 -473
rect 519 -507 587 -473
rect 677 -507 745 -473
rect 835 -507 903 -473
rect 993 -507 1061 -473
rect 1151 -507 1219 -473
rect 1309 -507 1377 -473
rect 1467 -507 1535 -473
rect 1625 -507 1693 -473
rect 1783 -507 1851 -473
rect 1941 -507 2009 -473
rect 2099 -507 2167 -473
rect -2229 -742 -2195 -566
rect -2071 -742 -2037 -566
rect -1913 -742 -1879 -566
rect -1755 -742 -1721 -566
rect -1597 -742 -1563 -566
rect -1439 -742 -1405 -566
rect -1281 -742 -1247 -566
rect -1123 -742 -1089 -566
rect -965 -742 -931 -566
rect -807 -742 -773 -566
rect -649 -742 -615 -566
rect -491 -742 -457 -566
rect -333 -742 -299 -566
rect -175 -742 -141 -566
rect -17 -742 17 -566
rect 141 -742 175 -566
rect 299 -742 333 -566
rect 457 -742 491 -566
rect 615 -742 649 -566
rect 773 -742 807 -566
rect 931 -742 965 -566
rect 1089 -742 1123 -566
rect 1247 -742 1281 -566
rect 1405 -742 1439 -566
rect 1563 -742 1597 -566
rect 1721 -742 1755 -566
rect 1879 -742 1913 -566
rect 2037 -742 2071 -566
rect 2195 -742 2229 -566
rect -2167 -835 -2099 -801
rect -2009 -835 -1941 -801
rect -1851 -835 -1783 -801
rect -1693 -835 -1625 -801
rect -1535 -835 -1467 -801
rect -1377 -835 -1309 -801
rect -1219 -835 -1151 -801
rect -1061 -835 -993 -801
rect -903 -835 -835 -801
rect -745 -835 -677 -801
rect -587 -835 -519 -801
rect -429 -835 -361 -801
rect -271 -835 -203 -801
rect -113 -835 -45 -801
rect 45 -835 113 -801
rect 203 -835 271 -801
rect 361 -835 429 -801
rect 519 -835 587 -801
rect 677 -835 745 -801
rect 835 -835 903 -801
rect 993 -835 1061 -801
rect 1151 -835 1219 -801
rect 1309 -835 1377 -801
rect 1467 -835 1535 -801
rect 1625 -835 1693 -801
rect 1783 -835 1851 -801
rect 1941 -835 2009 -801
rect 2099 -835 2167 -801
rect -2167 -943 -2099 -909
rect -2009 -943 -1941 -909
rect -1851 -943 -1783 -909
rect -1693 -943 -1625 -909
rect -1535 -943 -1467 -909
rect -1377 -943 -1309 -909
rect -1219 -943 -1151 -909
rect -1061 -943 -993 -909
rect -903 -943 -835 -909
rect -745 -943 -677 -909
rect -587 -943 -519 -909
rect -429 -943 -361 -909
rect -271 -943 -203 -909
rect -113 -943 -45 -909
rect 45 -943 113 -909
rect 203 -943 271 -909
rect 361 -943 429 -909
rect 519 -943 587 -909
rect 677 -943 745 -909
rect 835 -943 903 -909
rect 993 -943 1061 -909
rect 1151 -943 1219 -909
rect 1309 -943 1377 -909
rect 1467 -943 1535 -909
rect 1625 -943 1693 -909
rect 1783 -943 1851 -909
rect 1941 -943 2009 -909
rect 2099 -943 2167 -909
rect -2229 -1178 -2195 -1002
rect -2071 -1178 -2037 -1002
rect -1913 -1178 -1879 -1002
rect -1755 -1178 -1721 -1002
rect -1597 -1178 -1563 -1002
rect -1439 -1178 -1405 -1002
rect -1281 -1178 -1247 -1002
rect -1123 -1178 -1089 -1002
rect -965 -1178 -931 -1002
rect -807 -1178 -773 -1002
rect -649 -1178 -615 -1002
rect -491 -1178 -457 -1002
rect -333 -1178 -299 -1002
rect -175 -1178 -141 -1002
rect -17 -1178 17 -1002
rect 141 -1178 175 -1002
rect 299 -1178 333 -1002
rect 457 -1178 491 -1002
rect 615 -1178 649 -1002
rect 773 -1178 807 -1002
rect 931 -1178 965 -1002
rect 1089 -1178 1123 -1002
rect 1247 -1178 1281 -1002
rect 1405 -1178 1439 -1002
rect 1563 -1178 1597 -1002
rect 1721 -1178 1755 -1002
rect 1879 -1178 1913 -1002
rect 2037 -1178 2071 -1002
rect 2195 -1178 2229 -1002
rect -2167 -1271 -2099 -1237
rect -2009 -1271 -1941 -1237
rect -1851 -1271 -1783 -1237
rect -1693 -1271 -1625 -1237
rect -1535 -1271 -1467 -1237
rect -1377 -1271 -1309 -1237
rect -1219 -1271 -1151 -1237
rect -1061 -1271 -993 -1237
rect -903 -1271 -835 -1237
rect -745 -1271 -677 -1237
rect -587 -1271 -519 -1237
rect -429 -1271 -361 -1237
rect -271 -1271 -203 -1237
rect -113 -1271 -45 -1237
rect 45 -1271 113 -1237
rect 203 -1271 271 -1237
rect 361 -1271 429 -1237
rect 519 -1271 587 -1237
rect 677 -1271 745 -1237
rect 835 -1271 903 -1237
rect 993 -1271 1061 -1237
rect 1151 -1271 1219 -1237
rect 1309 -1271 1377 -1237
rect 1467 -1271 1535 -1237
rect 1625 -1271 1693 -1237
rect 1783 -1271 1851 -1237
rect 1941 -1271 2009 -1237
rect 2099 -1271 2167 -1237
rect -2167 -1379 -2099 -1345
rect -2009 -1379 -1941 -1345
rect -1851 -1379 -1783 -1345
rect -1693 -1379 -1625 -1345
rect -1535 -1379 -1467 -1345
rect -1377 -1379 -1309 -1345
rect -1219 -1379 -1151 -1345
rect -1061 -1379 -993 -1345
rect -903 -1379 -835 -1345
rect -745 -1379 -677 -1345
rect -587 -1379 -519 -1345
rect -429 -1379 -361 -1345
rect -271 -1379 -203 -1345
rect -113 -1379 -45 -1345
rect 45 -1379 113 -1345
rect 203 -1379 271 -1345
rect 361 -1379 429 -1345
rect 519 -1379 587 -1345
rect 677 -1379 745 -1345
rect 835 -1379 903 -1345
rect 993 -1379 1061 -1345
rect 1151 -1379 1219 -1345
rect 1309 -1379 1377 -1345
rect 1467 -1379 1535 -1345
rect 1625 -1379 1693 -1345
rect 1783 -1379 1851 -1345
rect 1941 -1379 2009 -1345
rect 2099 -1379 2167 -1345
rect -2229 -1614 -2195 -1438
rect -2071 -1614 -2037 -1438
rect -1913 -1614 -1879 -1438
rect -1755 -1614 -1721 -1438
rect -1597 -1614 -1563 -1438
rect -1439 -1614 -1405 -1438
rect -1281 -1614 -1247 -1438
rect -1123 -1614 -1089 -1438
rect -965 -1614 -931 -1438
rect -807 -1614 -773 -1438
rect -649 -1614 -615 -1438
rect -491 -1614 -457 -1438
rect -333 -1614 -299 -1438
rect -175 -1614 -141 -1438
rect -17 -1614 17 -1438
rect 141 -1614 175 -1438
rect 299 -1614 333 -1438
rect 457 -1614 491 -1438
rect 615 -1614 649 -1438
rect 773 -1614 807 -1438
rect 931 -1614 965 -1438
rect 1089 -1614 1123 -1438
rect 1247 -1614 1281 -1438
rect 1405 -1614 1439 -1438
rect 1563 -1614 1597 -1438
rect 1721 -1614 1755 -1438
rect 1879 -1614 1913 -1438
rect 2037 -1614 2071 -1438
rect 2195 -1614 2229 -1438
rect -2167 -1707 -2099 -1673
rect -2009 -1707 -1941 -1673
rect -1851 -1707 -1783 -1673
rect -1693 -1707 -1625 -1673
rect -1535 -1707 -1467 -1673
rect -1377 -1707 -1309 -1673
rect -1219 -1707 -1151 -1673
rect -1061 -1707 -993 -1673
rect -903 -1707 -835 -1673
rect -745 -1707 -677 -1673
rect -587 -1707 -519 -1673
rect -429 -1707 -361 -1673
rect -271 -1707 -203 -1673
rect -113 -1707 -45 -1673
rect 45 -1707 113 -1673
rect 203 -1707 271 -1673
rect 361 -1707 429 -1673
rect 519 -1707 587 -1673
rect 677 -1707 745 -1673
rect 835 -1707 903 -1673
rect 993 -1707 1061 -1673
rect 1151 -1707 1219 -1673
rect 1309 -1707 1377 -1673
rect 1467 -1707 1535 -1673
rect 1625 -1707 1693 -1673
rect 1783 -1707 1851 -1673
rect 1941 -1707 2009 -1673
rect 2099 -1707 2167 -1673
rect -2167 -1815 -2099 -1781
rect -2009 -1815 -1941 -1781
rect -1851 -1815 -1783 -1781
rect -1693 -1815 -1625 -1781
rect -1535 -1815 -1467 -1781
rect -1377 -1815 -1309 -1781
rect -1219 -1815 -1151 -1781
rect -1061 -1815 -993 -1781
rect -903 -1815 -835 -1781
rect -745 -1815 -677 -1781
rect -587 -1815 -519 -1781
rect -429 -1815 -361 -1781
rect -271 -1815 -203 -1781
rect -113 -1815 -45 -1781
rect 45 -1815 113 -1781
rect 203 -1815 271 -1781
rect 361 -1815 429 -1781
rect 519 -1815 587 -1781
rect 677 -1815 745 -1781
rect 835 -1815 903 -1781
rect 993 -1815 1061 -1781
rect 1151 -1815 1219 -1781
rect 1309 -1815 1377 -1781
rect 1467 -1815 1535 -1781
rect 1625 -1815 1693 -1781
rect 1783 -1815 1851 -1781
rect 1941 -1815 2009 -1781
rect 2099 -1815 2167 -1781
rect -2229 -2050 -2195 -1874
rect -2071 -2050 -2037 -1874
rect -1913 -2050 -1879 -1874
rect -1755 -2050 -1721 -1874
rect -1597 -2050 -1563 -1874
rect -1439 -2050 -1405 -1874
rect -1281 -2050 -1247 -1874
rect -1123 -2050 -1089 -1874
rect -965 -2050 -931 -1874
rect -807 -2050 -773 -1874
rect -649 -2050 -615 -1874
rect -491 -2050 -457 -1874
rect -333 -2050 -299 -1874
rect -175 -2050 -141 -1874
rect -17 -2050 17 -1874
rect 141 -2050 175 -1874
rect 299 -2050 333 -1874
rect 457 -2050 491 -1874
rect 615 -2050 649 -1874
rect 773 -2050 807 -1874
rect 931 -2050 965 -1874
rect 1089 -2050 1123 -1874
rect 1247 -2050 1281 -1874
rect 1405 -2050 1439 -1874
rect 1563 -2050 1597 -1874
rect 1721 -2050 1755 -1874
rect 1879 -2050 1913 -1874
rect 2037 -2050 2071 -1874
rect 2195 -2050 2229 -1874
rect -2167 -2143 -2099 -2109
rect -2009 -2143 -1941 -2109
rect -1851 -2143 -1783 -2109
rect -1693 -2143 -1625 -2109
rect -1535 -2143 -1467 -2109
rect -1377 -2143 -1309 -2109
rect -1219 -2143 -1151 -2109
rect -1061 -2143 -993 -2109
rect -903 -2143 -835 -2109
rect -745 -2143 -677 -2109
rect -587 -2143 -519 -2109
rect -429 -2143 -361 -2109
rect -271 -2143 -203 -2109
rect -113 -2143 -45 -2109
rect 45 -2143 113 -2109
rect 203 -2143 271 -2109
rect 361 -2143 429 -2109
rect 519 -2143 587 -2109
rect 677 -2143 745 -2109
rect 835 -2143 903 -2109
rect 993 -2143 1061 -2109
rect 1151 -2143 1219 -2109
rect 1309 -2143 1377 -2109
rect 1467 -2143 1535 -2109
rect 1625 -2143 1693 -2109
rect 1783 -2143 1851 -2109
rect 1941 -2143 2009 -2109
rect 2099 -2143 2167 -2109
<< metal1 >>
rect -2179 2143 -2087 2149
rect -2179 2109 -2167 2143
rect -2099 2109 -2087 2143
rect -2179 2103 -2087 2109
rect -2021 2143 -1929 2149
rect -2021 2109 -2009 2143
rect -1941 2109 -1929 2143
rect -2021 2103 -1929 2109
rect -1863 2143 -1771 2149
rect -1863 2109 -1851 2143
rect -1783 2109 -1771 2143
rect -1863 2103 -1771 2109
rect -1705 2143 -1613 2149
rect -1705 2109 -1693 2143
rect -1625 2109 -1613 2143
rect -1705 2103 -1613 2109
rect -1547 2143 -1455 2149
rect -1547 2109 -1535 2143
rect -1467 2109 -1455 2143
rect -1547 2103 -1455 2109
rect -1389 2143 -1297 2149
rect -1389 2109 -1377 2143
rect -1309 2109 -1297 2143
rect -1389 2103 -1297 2109
rect -1231 2143 -1139 2149
rect -1231 2109 -1219 2143
rect -1151 2109 -1139 2143
rect -1231 2103 -1139 2109
rect -1073 2143 -981 2149
rect -1073 2109 -1061 2143
rect -993 2109 -981 2143
rect -1073 2103 -981 2109
rect -915 2143 -823 2149
rect -915 2109 -903 2143
rect -835 2109 -823 2143
rect -915 2103 -823 2109
rect -757 2143 -665 2149
rect -757 2109 -745 2143
rect -677 2109 -665 2143
rect -757 2103 -665 2109
rect -599 2143 -507 2149
rect -599 2109 -587 2143
rect -519 2109 -507 2143
rect -599 2103 -507 2109
rect -441 2143 -349 2149
rect -441 2109 -429 2143
rect -361 2109 -349 2143
rect -441 2103 -349 2109
rect -283 2143 -191 2149
rect -283 2109 -271 2143
rect -203 2109 -191 2143
rect -283 2103 -191 2109
rect -125 2143 -33 2149
rect -125 2109 -113 2143
rect -45 2109 -33 2143
rect -125 2103 -33 2109
rect 33 2143 125 2149
rect 33 2109 45 2143
rect 113 2109 125 2143
rect 33 2103 125 2109
rect 191 2143 283 2149
rect 191 2109 203 2143
rect 271 2109 283 2143
rect 191 2103 283 2109
rect 349 2143 441 2149
rect 349 2109 361 2143
rect 429 2109 441 2143
rect 349 2103 441 2109
rect 507 2143 599 2149
rect 507 2109 519 2143
rect 587 2109 599 2143
rect 507 2103 599 2109
rect 665 2143 757 2149
rect 665 2109 677 2143
rect 745 2109 757 2143
rect 665 2103 757 2109
rect 823 2143 915 2149
rect 823 2109 835 2143
rect 903 2109 915 2143
rect 823 2103 915 2109
rect 981 2143 1073 2149
rect 981 2109 993 2143
rect 1061 2109 1073 2143
rect 981 2103 1073 2109
rect 1139 2143 1231 2149
rect 1139 2109 1151 2143
rect 1219 2109 1231 2143
rect 1139 2103 1231 2109
rect 1297 2143 1389 2149
rect 1297 2109 1309 2143
rect 1377 2109 1389 2143
rect 1297 2103 1389 2109
rect 1455 2143 1547 2149
rect 1455 2109 1467 2143
rect 1535 2109 1547 2143
rect 1455 2103 1547 2109
rect 1613 2143 1705 2149
rect 1613 2109 1625 2143
rect 1693 2109 1705 2143
rect 1613 2103 1705 2109
rect 1771 2143 1863 2149
rect 1771 2109 1783 2143
rect 1851 2109 1863 2143
rect 1771 2103 1863 2109
rect 1929 2143 2021 2149
rect 1929 2109 1941 2143
rect 2009 2109 2021 2143
rect 1929 2103 2021 2109
rect 2087 2143 2179 2149
rect 2087 2109 2099 2143
rect 2167 2109 2179 2143
rect 2087 2103 2179 2109
rect -2235 2050 -2189 2062
rect -2235 1874 -2229 2050
rect -2195 1874 -2189 2050
rect -2235 1862 -2189 1874
rect -2077 2050 -2031 2062
rect -2077 1874 -2071 2050
rect -2037 1874 -2031 2050
rect -2077 1862 -2031 1874
rect -1919 2050 -1873 2062
rect -1919 1874 -1913 2050
rect -1879 1874 -1873 2050
rect -1919 1862 -1873 1874
rect -1761 2050 -1715 2062
rect -1761 1874 -1755 2050
rect -1721 1874 -1715 2050
rect -1761 1862 -1715 1874
rect -1603 2050 -1557 2062
rect -1603 1874 -1597 2050
rect -1563 1874 -1557 2050
rect -1603 1862 -1557 1874
rect -1445 2050 -1399 2062
rect -1445 1874 -1439 2050
rect -1405 1874 -1399 2050
rect -1445 1862 -1399 1874
rect -1287 2050 -1241 2062
rect -1287 1874 -1281 2050
rect -1247 1874 -1241 2050
rect -1287 1862 -1241 1874
rect -1129 2050 -1083 2062
rect -1129 1874 -1123 2050
rect -1089 1874 -1083 2050
rect -1129 1862 -1083 1874
rect -971 2050 -925 2062
rect -971 1874 -965 2050
rect -931 1874 -925 2050
rect -971 1862 -925 1874
rect -813 2050 -767 2062
rect -813 1874 -807 2050
rect -773 1874 -767 2050
rect -813 1862 -767 1874
rect -655 2050 -609 2062
rect -655 1874 -649 2050
rect -615 1874 -609 2050
rect -655 1862 -609 1874
rect -497 2050 -451 2062
rect -497 1874 -491 2050
rect -457 1874 -451 2050
rect -497 1862 -451 1874
rect -339 2050 -293 2062
rect -339 1874 -333 2050
rect -299 1874 -293 2050
rect -339 1862 -293 1874
rect -181 2050 -135 2062
rect -181 1874 -175 2050
rect -141 1874 -135 2050
rect -181 1862 -135 1874
rect -23 2050 23 2062
rect -23 1874 -17 2050
rect 17 1874 23 2050
rect -23 1862 23 1874
rect 135 2050 181 2062
rect 135 1874 141 2050
rect 175 1874 181 2050
rect 135 1862 181 1874
rect 293 2050 339 2062
rect 293 1874 299 2050
rect 333 1874 339 2050
rect 293 1862 339 1874
rect 451 2050 497 2062
rect 451 1874 457 2050
rect 491 1874 497 2050
rect 451 1862 497 1874
rect 609 2050 655 2062
rect 609 1874 615 2050
rect 649 1874 655 2050
rect 609 1862 655 1874
rect 767 2050 813 2062
rect 767 1874 773 2050
rect 807 1874 813 2050
rect 767 1862 813 1874
rect 925 2050 971 2062
rect 925 1874 931 2050
rect 965 1874 971 2050
rect 925 1862 971 1874
rect 1083 2050 1129 2062
rect 1083 1874 1089 2050
rect 1123 1874 1129 2050
rect 1083 1862 1129 1874
rect 1241 2050 1287 2062
rect 1241 1874 1247 2050
rect 1281 1874 1287 2050
rect 1241 1862 1287 1874
rect 1399 2050 1445 2062
rect 1399 1874 1405 2050
rect 1439 1874 1445 2050
rect 1399 1862 1445 1874
rect 1557 2050 1603 2062
rect 1557 1874 1563 2050
rect 1597 1874 1603 2050
rect 1557 1862 1603 1874
rect 1715 2050 1761 2062
rect 1715 1874 1721 2050
rect 1755 1874 1761 2050
rect 1715 1862 1761 1874
rect 1873 2050 1919 2062
rect 1873 1874 1879 2050
rect 1913 1874 1919 2050
rect 1873 1862 1919 1874
rect 2031 2050 2077 2062
rect 2031 1874 2037 2050
rect 2071 1874 2077 2050
rect 2031 1862 2077 1874
rect 2189 2050 2235 2062
rect 2189 1874 2195 2050
rect 2229 1874 2235 2050
rect 2189 1862 2235 1874
rect -2179 1815 -2087 1821
rect -2179 1781 -2167 1815
rect -2099 1781 -2087 1815
rect -2179 1775 -2087 1781
rect -2021 1815 -1929 1821
rect -2021 1781 -2009 1815
rect -1941 1781 -1929 1815
rect -2021 1775 -1929 1781
rect -1863 1815 -1771 1821
rect -1863 1781 -1851 1815
rect -1783 1781 -1771 1815
rect -1863 1775 -1771 1781
rect -1705 1815 -1613 1821
rect -1705 1781 -1693 1815
rect -1625 1781 -1613 1815
rect -1705 1775 -1613 1781
rect -1547 1815 -1455 1821
rect -1547 1781 -1535 1815
rect -1467 1781 -1455 1815
rect -1547 1775 -1455 1781
rect -1389 1815 -1297 1821
rect -1389 1781 -1377 1815
rect -1309 1781 -1297 1815
rect -1389 1775 -1297 1781
rect -1231 1815 -1139 1821
rect -1231 1781 -1219 1815
rect -1151 1781 -1139 1815
rect -1231 1775 -1139 1781
rect -1073 1815 -981 1821
rect -1073 1781 -1061 1815
rect -993 1781 -981 1815
rect -1073 1775 -981 1781
rect -915 1815 -823 1821
rect -915 1781 -903 1815
rect -835 1781 -823 1815
rect -915 1775 -823 1781
rect -757 1815 -665 1821
rect -757 1781 -745 1815
rect -677 1781 -665 1815
rect -757 1775 -665 1781
rect -599 1815 -507 1821
rect -599 1781 -587 1815
rect -519 1781 -507 1815
rect -599 1775 -507 1781
rect -441 1815 -349 1821
rect -441 1781 -429 1815
rect -361 1781 -349 1815
rect -441 1775 -349 1781
rect -283 1815 -191 1821
rect -283 1781 -271 1815
rect -203 1781 -191 1815
rect -283 1775 -191 1781
rect -125 1815 -33 1821
rect -125 1781 -113 1815
rect -45 1781 -33 1815
rect -125 1775 -33 1781
rect 33 1815 125 1821
rect 33 1781 45 1815
rect 113 1781 125 1815
rect 33 1775 125 1781
rect 191 1815 283 1821
rect 191 1781 203 1815
rect 271 1781 283 1815
rect 191 1775 283 1781
rect 349 1815 441 1821
rect 349 1781 361 1815
rect 429 1781 441 1815
rect 349 1775 441 1781
rect 507 1815 599 1821
rect 507 1781 519 1815
rect 587 1781 599 1815
rect 507 1775 599 1781
rect 665 1815 757 1821
rect 665 1781 677 1815
rect 745 1781 757 1815
rect 665 1775 757 1781
rect 823 1815 915 1821
rect 823 1781 835 1815
rect 903 1781 915 1815
rect 823 1775 915 1781
rect 981 1815 1073 1821
rect 981 1781 993 1815
rect 1061 1781 1073 1815
rect 981 1775 1073 1781
rect 1139 1815 1231 1821
rect 1139 1781 1151 1815
rect 1219 1781 1231 1815
rect 1139 1775 1231 1781
rect 1297 1815 1389 1821
rect 1297 1781 1309 1815
rect 1377 1781 1389 1815
rect 1297 1775 1389 1781
rect 1455 1815 1547 1821
rect 1455 1781 1467 1815
rect 1535 1781 1547 1815
rect 1455 1775 1547 1781
rect 1613 1815 1705 1821
rect 1613 1781 1625 1815
rect 1693 1781 1705 1815
rect 1613 1775 1705 1781
rect 1771 1815 1863 1821
rect 1771 1781 1783 1815
rect 1851 1781 1863 1815
rect 1771 1775 1863 1781
rect 1929 1815 2021 1821
rect 1929 1781 1941 1815
rect 2009 1781 2021 1815
rect 1929 1775 2021 1781
rect 2087 1815 2179 1821
rect 2087 1781 2099 1815
rect 2167 1781 2179 1815
rect 2087 1775 2179 1781
rect -2179 1707 -2087 1713
rect -2179 1673 -2167 1707
rect -2099 1673 -2087 1707
rect -2179 1667 -2087 1673
rect -2021 1707 -1929 1713
rect -2021 1673 -2009 1707
rect -1941 1673 -1929 1707
rect -2021 1667 -1929 1673
rect -1863 1707 -1771 1713
rect -1863 1673 -1851 1707
rect -1783 1673 -1771 1707
rect -1863 1667 -1771 1673
rect -1705 1707 -1613 1713
rect -1705 1673 -1693 1707
rect -1625 1673 -1613 1707
rect -1705 1667 -1613 1673
rect -1547 1707 -1455 1713
rect -1547 1673 -1535 1707
rect -1467 1673 -1455 1707
rect -1547 1667 -1455 1673
rect -1389 1707 -1297 1713
rect -1389 1673 -1377 1707
rect -1309 1673 -1297 1707
rect -1389 1667 -1297 1673
rect -1231 1707 -1139 1713
rect -1231 1673 -1219 1707
rect -1151 1673 -1139 1707
rect -1231 1667 -1139 1673
rect -1073 1707 -981 1713
rect -1073 1673 -1061 1707
rect -993 1673 -981 1707
rect -1073 1667 -981 1673
rect -915 1707 -823 1713
rect -915 1673 -903 1707
rect -835 1673 -823 1707
rect -915 1667 -823 1673
rect -757 1707 -665 1713
rect -757 1673 -745 1707
rect -677 1673 -665 1707
rect -757 1667 -665 1673
rect -599 1707 -507 1713
rect -599 1673 -587 1707
rect -519 1673 -507 1707
rect -599 1667 -507 1673
rect -441 1707 -349 1713
rect -441 1673 -429 1707
rect -361 1673 -349 1707
rect -441 1667 -349 1673
rect -283 1707 -191 1713
rect -283 1673 -271 1707
rect -203 1673 -191 1707
rect -283 1667 -191 1673
rect -125 1707 -33 1713
rect -125 1673 -113 1707
rect -45 1673 -33 1707
rect -125 1667 -33 1673
rect 33 1707 125 1713
rect 33 1673 45 1707
rect 113 1673 125 1707
rect 33 1667 125 1673
rect 191 1707 283 1713
rect 191 1673 203 1707
rect 271 1673 283 1707
rect 191 1667 283 1673
rect 349 1707 441 1713
rect 349 1673 361 1707
rect 429 1673 441 1707
rect 349 1667 441 1673
rect 507 1707 599 1713
rect 507 1673 519 1707
rect 587 1673 599 1707
rect 507 1667 599 1673
rect 665 1707 757 1713
rect 665 1673 677 1707
rect 745 1673 757 1707
rect 665 1667 757 1673
rect 823 1707 915 1713
rect 823 1673 835 1707
rect 903 1673 915 1707
rect 823 1667 915 1673
rect 981 1707 1073 1713
rect 981 1673 993 1707
rect 1061 1673 1073 1707
rect 981 1667 1073 1673
rect 1139 1707 1231 1713
rect 1139 1673 1151 1707
rect 1219 1673 1231 1707
rect 1139 1667 1231 1673
rect 1297 1707 1389 1713
rect 1297 1673 1309 1707
rect 1377 1673 1389 1707
rect 1297 1667 1389 1673
rect 1455 1707 1547 1713
rect 1455 1673 1467 1707
rect 1535 1673 1547 1707
rect 1455 1667 1547 1673
rect 1613 1707 1705 1713
rect 1613 1673 1625 1707
rect 1693 1673 1705 1707
rect 1613 1667 1705 1673
rect 1771 1707 1863 1713
rect 1771 1673 1783 1707
rect 1851 1673 1863 1707
rect 1771 1667 1863 1673
rect 1929 1707 2021 1713
rect 1929 1673 1941 1707
rect 2009 1673 2021 1707
rect 1929 1667 2021 1673
rect 2087 1707 2179 1713
rect 2087 1673 2099 1707
rect 2167 1673 2179 1707
rect 2087 1667 2179 1673
rect -2235 1614 -2189 1626
rect -2235 1438 -2229 1614
rect -2195 1438 -2189 1614
rect -2235 1426 -2189 1438
rect -2077 1614 -2031 1626
rect -2077 1438 -2071 1614
rect -2037 1438 -2031 1614
rect -2077 1426 -2031 1438
rect -1919 1614 -1873 1626
rect -1919 1438 -1913 1614
rect -1879 1438 -1873 1614
rect -1919 1426 -1873 1438
rect -1761 1614 -1715 1626
rect -1761 1438 -1755 1614
rect -1721 1438 -1715 1614
rect -1761 1426 -1715 1438
rect -1603 1614 -1557 1626
rect -1603 1438 -1597 1614
rect -1563 1438 -1557 1614
rect -1603 1426 -1557 1438
rect -1445 1614 -1399 1626
rect -1445 1438 -1439 1614
rect -1405 1438 -1399 1614
rect -1445 1426 -1399 1438
rect -1287 1614 -1241 1626
rect -1287 1438 -1281 1614
rect -1247 1438 -1241 1614
rect -1287 1426 -1241 1438
rect -1129 1614 -1083 1626
rect -1129 1438 -1123 1614
rect -1089 1438 -1083 1614
rect -1129 1426 -1083 1438
rect -971 1614 -925 1626
rect -971 1438 -965 1614
rect -931 1438 -925 1614
rect -971 1426 -925 1438
rect -813 1614 -767 1626
rect -813 1438 -807 1614
rect -773 1438 -767 1614
rect -813 1426 -767 1438
rect -655 1614 -609 1626
rect -655 1438 -649 1614
rect -615 1438 -609 1614
rect -655 1426 -609 1438
rect -497 1614 -451 1626
rect -497 1438 -491 1614
rect -457 1438 -451 1614
rect -497 1426 -451 1438
rect -339 1614 -293 1626
rect -339 1438 -333 1614
rect -299 1438 -293 1614
rect -339 1426 -293 1438
rect -181 1614 -135 1626
rect -181 1438 -175 1614
rect -141 1438 -135 1614
rect -181 1426 -135 1438
rect -23 1614 23 1626
rect -23 1438 -17 1614
rect 17 1438 23 1614
rect -23 1426 23 1438
rect 135 1614 181 1626
rect 135 1438 141 1614
rect 175 1438 181 1614
rect 135 1426 181 1438
rect 293 1614 339 1626
rect 293 1438 299 1614
rect 333 1438 339 1614
rect 293 1426 339 1438
rect 451 1614 497 1626
rect 451 1438 457 1614
rect 491 1438 497 1614
rect 451 1426 497 1438
rect 609 1614 655 1626
rect 609 1438 615 1614
rect 649 1438 655 1614
rect 609 1426 655 1438
rect 767 1614 813 1626
rect 767 1438 773 1614
rect 807 1438 813 1614
rect 767 1426 813 1438
rect 925 1614 971 1626
rect 925 1438 931 1614
rect 965 1438 971 1614
rect 925 1426 971 1438
rect 1083 1614 1129 1626
rect 1083 1438 1089 1614
rect 1123 1438 1129 1614
rect 1083 1426 1129 1438
rect 1241 1614 1287 1626
rect 1241 1438 1247 1614
rect 1281 1438 1287 1614
rect 1241 1426 1287 1438
rect 1399 1614 1445 1626
rect 1399 1438 1405 1614
rect 1439 1438 1445 1614
rect 1399 1426 1445 1438
rect 1557 1614 1603 1626
rect 1557 1438 1563 1614
rect 1597 1438 1603 1614
rect 1557 1426 1603 1438
rect 1715 1614 1761 1626
rect 1715 1438 1721 1614
rect 1755 1438 1761 1614
rect 1715 1426 1761 1438
rect 1873 1614 1919 1626
rect 1873 1438 1879 1614
rect 1913 1438 1919 1614
rect 1873 1426 1919 1438
rect 2031 1614 2077 1626
rect 2031 1438 2037 1614
rect 2071 1438 2077 1614
rect 2031 1426 2077 1438
rect 2189 1614 2235 1626
rect 2189 1438 2195 1614
rect 2229 1438 2235 1614
rect 2189 1426 2235 1438
rect -2179 1379 -2087 1385
rect -2179 1345 -2167 1379
rect -2099 1345 -2087 1379
rect -2179 1339 -2087 1345
rect -2021 1379 -1929 1385
rect -2021 1345 -2009 1379
rect -1941 1345 -1929 1379
rect -2021 1339 -1929 1345
rect -1863 1379 -1771 1385
rect -1863 1345 -1851 1379
rect -1783 1345 -1771 1379
rect -1863 1339 -1771 1345
rect -1705 1379 -1613 1385
rect -1705 1345 -1693 1379
rect -1625 1345 -1613 1379
rect -1705 1339 -1613 1345
rect -1547 1379 -1455 1385
rect -1547 1345 -1535 1379
rect -1467 1345 -1455 1379
rect -1547 1339 -1455 1345
rect -1389 1379 -1297 1385
rect -1389 1345 -1377 1379
rect -1309 1345 -1297 1379
rect -1389 1339 -1297 1345
rect -1231 1379 -1139 1385
rect -1231 1345 -1219 1379
rect -1151 1345 -1139 1379
rect -1231 1339 -1139 1345
rect -1073 1379 -981 1385
rect -1073 1345 -1061 1379
rect -993 1345 -981 1379
rect -1073 1339 -981 1345
rect -915 1379 -823 1385
rect -915 1345 -903 1379
rect -835 1345 -823 1379
rect -915 1339 -823 1345
rect -757 1379 -665 1385
rect -757 1345 -745 1379
rect -677 1345 -665 1379
rect -757 1339 -665 1345
rect -599 1379 -507 1385
rect -599 1345 -587 1379
rect -519 1345 -507 1379
rect -599 1339 -507 1345
rect -441 1379 -349 1385
rect -441 1345 -429 1379
rect -361 1345 -349 1379
rect -441 1339 -349 1345
rect -283 1379 -191 1385
rect -283 1345 -271 1379
rect -203 1345 -191 1379
rect -283 1339 -191 1345
rect -125 1379 -33 1385
rect -125 1345 -113 1379
rect -45 1345 -33 1379
rect -125 1339 -33 1345
rect 33 1379 125 1385
rect 33 1345 45 1379
rect 113 1345 125 1379
rect 33 1339 125 1345
rect 191 1379 283 1385
rect 191 1345 203 1379
rect 271 1345 283 1379
rect 191 1339 283 1345
rect 349 1379 441 1385
rect 349 1345 361 1379
rect 429 1345 441 1379
rect 349 1339 441 1345
rect 507 1379 599 1385
rect 507 1345 519 1379
rect 587 1345 599 1379
rect 507 1339 599 1345
rect 665 1379 757 1385
rect 665 1345 677 1379
rect 745 1345 757 1379
rect 665 1339 757 1345
rect 823 1379 915 1385
rect 823 1345 835 1379
rect 903 1345 915 1379
rect 823 1339 915 1345
rect 981 1379 1073 1385
rect 981 1345 993 1379
rect 1061 1345 1073 1379
rect 981 1339 1073 1345
rect 1139 1379 1231 1385
rect 1139 1345 1151 1379
rect 1219 1345 1231 1379
rect 1139 1339 1231 1345
rect 1297 1379 1389 1385
rect 1297 1345 1309 1379
rect 1377 1345 1389 1379
rect 1297 1339 1389 1345
rect 1455 1379 1547 1385
rect 1455 1345 1467 1379
rect 1535 1345 1547 1379
rect 1455 1339 1547 1345
rect 1613 1379 1705 1385
rect 1613 1345 1625 1379
rect 1693 1345 1705 1379
rect 1613 1339 1705 1345
rect 1771 1379 1863 1385
rect 1771 1345 1783 1379
rect 1851 1345 1863 1379
rect 1771 1339 1863 1345
rect 1929 1379 2021 1385
rect 1929 1345 1941 1379
rect 2009 1345 2021 1379
rect 1929 1339 2021 1345
rect 2087 1379 2179 1385
rect 2087 1345 2099 1379
rect 2167 1345 2179 1379
rect 2087 1339 2179 1345
rect -2179 1271 -2087 1277
rect -2179 1237 -2167 1271
rect -2099 1237 -2087 1271
rect -2179 1231 -2087 1237
rect -2021 1271 -1929 1277
rect -2021 1237 -2009 1271
rect -1941 1237 -1929 1271
rect -2021 1231 -1929 1237
rect -1863 1271 -1771 1277
rect -1863 1237 -1851 1271
rect -1783 1237 -1771 1271
rect -1863 1231 -1771 1237
rect -1705 1271 -1613 1277
rect -1705 1237 -1693 1271
rect -1625 1237 -1613 1271
rect -1705 1231 -1613 1237
rect -1547 1271 -1455 1277
rect -1547 1237 -1535 1271
rect -1467 1237 -1455 1271
rect -1547 1231 -1455 1237
rect -1389 1271 -1297 1277
rect -1389 1237 -1377 1271
rect -1309 1237 -1297 1271
rect -1389 1231 -1297 1237
rect -1231 1271 -1139 1277
rect -1231 1237 -1219 1271
rect -1151 1237 -1139 1271
rect -1231 1231 -1139 1237
rect -1073 1271 -981 1277
rect -1073 1237 -1061 1271
rect -993 1237 -981 1271
rect -1073 1231 -981 1237
rect -915 1271 -823 1277
rect -915 1237 -903 1271
rect -835 1237 -823 1271
rect -915 1231 -823 1237
rect -757 1271 -665 1277
rect -757 1237 -745 1271
rect -677 1237 -665 1271
rect -757 1231 -665 1237
rect -599 1271 -507 1277
rect -599 1237 -587 1271
rect -519 1237 -507 1271
rect -599 1231 -507 1237
rect -441 1271 -349 1277
rect -441 1237 -429 1271
rect -361 1237 -349 1271
rect -441 1231 -349 1237
rect -283 1271 -191 1277
rect -283 1237 -271 1271
rect -203 1237 -191 1271
rect -283 1231 -191 1237
rect -125 1271 -33 1277
rect -125 1237 -113 1271
rect -45 1237 -33 1271
rect -125 1231 -33 1237
rect 33 1271 125 1277
rect 33 1237 45 1271
rect 113 1237 125 1271
rect 33 1231 125 1237
rect 191 1271 283 1277
rect 191 1237 203 1271
rect 271 1237 283 1271
rect 191 1231 283 1237
rect 349 1271 441 1277
rect 349 1237 361 1271
rect 429 1237 441 1271
rect 349 1231 441 1237
rect 507 1271 599 1277
rect 507 1237 519 1271
rect 587 1237 599 1271
rect 507 1231 599 1237
rect 665 1271 757 1277
rect 665 1237 677 1271
rect 745 1237 757 1271
rect 665 1231 757 1237
rect 823 1271 915 1277
rect 823 1237 835 1271
rect 903 1237 915 1271
rect 823 1231 915 1237
rect 981 1271 1073 1277
rect 981 1237 993 1271
rect 1061 1237 1073 1271
rect 981 1231 1073 1237
rect 1139 1271 1231 1277
rect 1139 1237 1151 1271
rect 1219 1237 1231 1271
rect 1139 1231 1231 1237
rect 1297 1271 1389 1277
rect 1297 1237 1309 1271
rect 1377 1237 1389 1271
rect 1297 1231 1389 1237
rect 1455 1271 1547 1277
rect 1455 1237 1467 1271
rect 1535 1237 1547 1271
rect 1455 1231 1547 1237
rect 1613 1271 1705 1277
rect 1613 1237 1625 1271
rect 1693 1237 1705 1271
rect 1613 1231 1705 1237
rect 1771 1271 1863 1277
rect 1771 1237 1783 1271
rect 1851 1237 1863 1271
rect 1771 1231 1863 1237
rect 1929 1271 2021 1277
rect 1929 1237 1941 1271
rect 2009 1237 2021 1271
rect 1929 1231 2021 1237
rect 2087 1271 2179 1277
rect 2087 1237 2099 1271
rect 2167 1237 2179 1271
rect 2087 1231 2179 1237
rect -2235 1178 -2189 1190
rect -2235 1002 -2229 1178
rect -2195 1002 -2189 1178
rect -2235 990 -2189 1002
rect -2077 1178 -2031 1190
rect -2077 1002 -2071 1178
rect -2037 1002 -2031 1178
rect -2077 990 -2031 1002
rect -1919 1178 -1873 1190
rect -1919 1002 -1913 1178
rect -1879 1002 -1873 1178
rect -1919 990 -1873 1002
rect -1761 1178 -1715 1190
rect -1761 1002 -1755 1178
rect -1721 1002 -1715 1178
rect -1761 990 -1715 1002
rect -1603 1178 -1557 1190
rect -1603 1002 -1597 1178
rect -1563 1002 -1557 1178
rect -1603 990 -1557 1002
rect -1445 1178 -1399 1190
rect -1445 1002 -1439 1178
rect -1405 1002 -1399 1178
rect -1445 990 -1399 1002
rect -1287 1178 -1241 1190
rect -1287 1002 -1281 1178
rect -1247 1002 -1241 1178
rect -1287 990 -1241 1002
rect -1129 1178 -1083 1190
rect -1129 1002 -1123 1178
rect -1089 1002 -1083 1178
rect -1129 990 -1083 1002
rect -971 1178 -925 1190
rect -971 1002 -965 1178
rect -931 1002 -925 1178
rect -971 990 -925 1002
rect -813 1178 -767 1190
rect -813 1002 -807 1178
rect -773 1002 -767 1178
rect -813 990 -767 1002
rect -655 1178 -609 1190
rect -655 1002 -649 1178
rect -615 1002 -609 1178
rect -655 990 -609 1002
rect -497 1178 -451 1190
rect -497 1002 -491 1178
rect -457 1002 -451 1178
rect -497 990 -451 1002
rect -339 1178 -293 1190
rect -339 1002 -333 1178
rect -299 1002 -293 1178
rect -339 990 -293 1002
rect -181 1178 -135 1190
rect -181 1002 -175 1178
rect -141 1002 -135 1178
rect -181 990 -135 1002
rect -23 1178 23 1190
rect -23 1002 -17 1178
rect 17 1002 23 1178
rect -23 990 23 1002
rect 135 1178 181 1190
rect 135 1002 141 1178
rect 175 1002 181 1178
rect 135 990 181 1002
rect 293 1178 339 1190
rect 293 1002 299 1178
rect 333 1002 339 1178
rect 293 990 339 1002
rect 451 1178 497 1190
rect 451 1002 457 1178
rect 491 1002 497 1178
rect 451 990 497 1002
rect 609 1178 655 1190
rect 609 1002 615 1178
rect 649 1002 655 1178
rect 609 990 655 1002
rect 767 1178 813 1190
rect 767 1002 773 1178
rect 807 1002 813 1178
rect 767 990 813 1002
rect 925 1178 971 1190
rect 925 1002 931 1178
rect 965 1002 971 1178
rect 925 990 971 1002
rect 1083 1178 1129 1190
rect 1083 1002 1089 1178
rect 1123 1002 1129 1178
rect 1083 990 1129 1002
rect 1241 1178 1287 1190
rect 1241 1002 1247 1178
rect 1281 1002 1287 1178
rect 1241 990 1287 1002
rect 1399 1178 1445 1190
rect 1399 1002 1405 1178
rect 1439 1002 1445 1178
rect 1399 990 1445 1002
rect 1557 1178 1603 1190
rect 1557 1002 1563 1178
rect 1597 1002 1603 1178
rect 1557 990 1603 1002
rect 1715 1178 1761 1190
rect 1715 1002 1721 1178
rect 1755 1002 1761 1178
rect 1715 990 1761 1002
rect 1873 1178 1919 1190
rect 1873 1002 1879 1178
rect 1913 1002 1919 1178
rect 1873 990 1919 1002
rect 2031 1178 2077 1190
rect 2031 1002 2037 1178
rect 2071 1002 2077 1178
rect 2031 990 2077 1002
rect 2189 1178 2235 1190
rect 2189 1002 2195 1178
rect 2229 1002 2235 1178
rect 2189 990 2235 1002
rect -2179 943 -2087 949
rect -2179 909 -2167 943
rect -2099 909 -2087 943
rect -2179 903 -2087 909
rect -2021 943 -1929 949
rect -2021 909 -2009 943
rect -1941 909 -1929 943
rect -2021 903 -1929 909
rect -1863 943 -1771 949
rect -1863 909 -1851 943
rect -1783 909 -1771 943
rect -1863 903 -1771 909
rect -1705 943 -1613 949
rect -1705 909 -1693 943
rect -1625 909 -1613 943
rect -1705 903 -1613 909
rect -1547 943 -1455 949
rect -1547 909 -1535 943
rect -1467 909 -1455 943
rect -1547 903 -1455 909
rect -1389 943 -1297 949
rect -1389 909 -1377 943
rect -1309 909 -1297 943
rect -1389 903 -1297 909
rect -1231 943 -1139 949
rect -1231 909 -1219 943
rect -1151 909 -1139 943
rect -1231 903 -1139 909
rect -1073 943 -981 949
rect -1073 909 -1061 943
rect -993 909 -981 943
rect -1073 903 -981 909
rect -915 943 -823 949
rect -915 909 -903 943
rect -835 909 -823 943
rect -915 903 -823 909
rect -757 943 -665 949
rect -757 909 -745 943
rect -677 909 -665 943
rect -757 903 -665 909
rect -599 943 -507 949
rect -599 909 -587 943
rect -519 909 -507 943
rect -599 903 -507 909
rect -441 943 -349 949
rect -441 909 -429 943
rect -361 909 -349 943
rect -441 903 -349 909
rect -283 943 -191 949
rect -283 909 -271 943
rect -203 909 -191 943
rect -283 903 -191 909
rect -125 943 -33 949
rect -125 909 -113 943
rect -45 909 -33 943
rect -125 903 -33 909
rect 33 943 125 949
rect 33 909 45 943
rect 113 909 125 943
rect 33 903 125 909
rect 191 943 283 949
rect 191 909 203 943
rect 271 909 283 943
rect 191 903 283 909
rect 349 943 441 949
rect 349 909 361 943
rect 429 909 441 943
rect 349 903 441 909
rect 507 943 599 949
rect 507 909 519 943
rect 587 909 599 943
rect 507 903 599 909
rect 665 943 757 949
rect 665 909 677 943
rect 745 909 757 943
rect 665 903 757 909
rect 823 943 915 949
rect 823 909 835 943
rect 903 909 915 943
rect 823 903 915 909
rect 981 943 1073 949
rect 981 909 993 943
rect 1061 909 1073 943
rect 981 903 1073 909
rect 1139 943 1231 949
rect 1139 909 1151 943
rect 1219 909 1231 943
rect 1139 903 1231 909
rect 1297 943 1389 949
rect 1297 909 1309 943
rect 1377 909 1389 943
rect 1297 903 1389 909
rect 1455 943 1547 949
rect 1455 909 1467 943
rect 1535 909 1547 943
rect 1455 903 1547 909
rect 1613 943 1705 949
rect 1613 909 1625 943
rect 1693 909 1705 943
rect 1613 903 1705 909
rect 1771 943 1863 949
rect 1771 909 1783 943
rect 1851 909 1863 943
rect 1771 903 1863 909
rect 1929 943 2021 949
rect 1929 909 1941 943
rect 2009 909 2021 943
rect 1929 903 2021 909
rect 2087 943 2179 949
rect 2087 909 2099 943
rect 2167 909 2179 943
rect 2087 903 2179 909
rect -2179 835 -2087 841
rect -2179 801 -2167 835
rect -2099 801 -2087 835
rect -2179 795 -2087 801
rect -2021 835 -1929 841
rect -2021 801 -2009 835
rect -1941 801 -1929 835
rect -2021 795 -1929 801
rect -1863 835 -1771 841
rect -1863 801 -1851 835
rect -1783 801 -1771 835
rect -1863 795 -1771 801
rect -1705 835 -1613 841
rect -1705 801 -1693 835
rect -1625 801 -1613 835
rect -1705 795 -1613 801
rect -1547 835 -1455 841
rect -1547 801 -1535 835
rect -1467 801 -1455 835
rect -1547 795 -1455 801
rect -1389 835 -1297 841
rect -1389 801 -1377 835
rect -1309 801 -1297 835
rect -1389 795 -1297 801
rect -1231 835 -1139 841
rect -1231 801 -1219 835
rect -1151 801 -1139 835
rect -1231 795 -1139 801
rect -1073 835 -981 841
rect -1073 801 -1061 835
rect -993 801 -981 835
rect -1073 795 -981 801
rect -915 835 -823 841
rect -915 801 -903 835
rect -835 801 -823 835
rect -915 795 -823 801
rect -757 835 -665 841
rect -757 801 -745 835
rect -677 801 -665 835
rect -757 795 -665 801
rect -599 835 -507 841
rect -599 801 -587 835
rect -519 801 -507 835
rect -599 795 -507 801
rect -441 835 -349 841
rect -441 801 -429 835
rect -361 801 -349 835
rect -441 795 -349 801
rect -283 835 -191 841
rect -283 801 -271 835
rect -203 801 -191 835
rect -283 795 -191 801
rect -125 835 -33 841
rect -125 801 -113 835
rect -45 801 -33 835
rect -125 795 -33 801
rect 33 835 125 841
rect 33 801 45 835
rect 113 801 125 835
rect 33 795 125 801
rect 191 835 283 841
rect 191 801 203 835
rect 271 801 283 835
rect 191 795 283 801
rect 349 835 441 841
rect 349 801 361 835
rect 429 801 441 835
rect 349 795 441 801
rect 507 835 599 841
rect 507 801 519 835
rect 587 801 599 835
rect 507 795 599 801
rect 665 835 757 841
rect 665 801 677 835
rect 745 801 757 835
rect 665 795 757 801
rect 823 835 915 841
rect 823 801 835 835
rect 903 801 915 835
rect 823 795 915 801
rect 981 835 1073 841
rect 981 801 993 835
rect 1061 801 1073 835
rect 981 795 1073 801
rect 1139 835 1231 841
rect 1139 801 1151 835
rect 1219 801 1231 835
rect 1139 795 1231 801
rect 1297 835 1389 841
rect 1297 801 1309 835
rect 1377 801 1389 835
rect 1297 795 1389 801
rect 1455 835 1547 841
rect 1455 801 1467 835
rect 1535 801 1547 835
rect 1455 795 1547 801
rect 1613 835 1705 841
rect 1613 801 1625 835
rect 1693 801 1705 835
rect 1613 795 1705 801
rect 1771 835 1863 841
rect 1771 801 1783 835
rect 1851 801 1863 835
rect 1771 795 1863 801
rect 1929 835 2021 841
rect 1929 801 1941 835
rect 2009 801 2021 835
rect 1929 795 2021 801
rect 2087 835 2179 841
rect 2087 801 2099 835
rect 2167 801 2179 835
rect 2087 795 2179 801
rect -2235 742 -2189 754
rect -2235 566 -2229 742
rect -2195 566 -2189 742
rect -2235 554 -2189 566
rect -2077 742 -2031 754
rect -2077 566 -2071 742
rect -2037 566 -2031 742
rect -2077 554 -2031 566
rect -1919 742 -1873 754
rect -1919 566 -1913 742
rect -1879 566 -1873 742
rect -1919 554 -1873 566
rect -1761 742 -1715 754
rect -1761 566 -1755 742
rect -1721 566 -1715 742
rect -1761 554 -1715 566
rect -1603 742 -1557 754
rect -1603 566 -1597 742
rect -1563 566 -1557 742
rect -1603 554 -1557 566
rect -1445 742 -1399 754
rect -1445 566 -1439 742
rect -1405 566 -1399 742
rect -1445 554 -1399 566
rect -1287 742 -1241 754
rect -1287 566 -1281 742
rect -1247 566 -1241 742
rect -1287 554 -1241 566
rect -1129 742 -1083 754
rect -1129 566 -1123 742
rect -1089 566 -1083 742
rect -1129 554 -1083 566
rect -971 742 -925 754
rect -971 566 -965 742
rect -931 566 -925 742
rect -971 554 -925 566
rect -813 742 -767 754
rect -813 566 -807 742
rect -773 566 -767 742
rect -813 554 -767 566
rect -655 742 -609 754
rect -655 566 -649 742
rect -615 566 -609 742
rect -655 554 -609 566
rect -497 742 -451 754
rect -497 566 -491 742
rect -457 566 -451 742
rect -497 554 -451 566
rect -339 742 -293 754
rect -339 566 -333 742
rect -299 566 -293 742
rect -339 554 -293 566
rect -181 742 -135 754
rect -181 566 -175 742
rect -141 566 -135 742
rect -181 554 -135 566
rect -23 742 23 754
rect -23 566 -17 742
rect 17 566 23 742
rect -23 554 23 566
rect 135 742 181 754
rect 135 566 141 742
rect 175 566 181 742
rect 135 554 181 566
rect 293 742 339 754
rect 293 566 299 742
rect 333 566 339 742
rect 293 554 339 566
rect 451 742 497 754
rect 451 566 457 742
rect 491 566 497 742
rect 451 554 497 566
rect 609 742 655 754
rect 609 566 615 742
rect 649 566 655 742
rect 609 554 655 566
rect 767 742 813 754
rect 767 566 773 742
rect 807 566 813 742
rect 767 554 813 566
rect 925 742 971 754
rect 925 566 931 742
rect 965 566 971 742
rect 925 554 971 566
rect 1083 742 1129 754
rect 1083 566 1089 742
rect 1123 566 1129 742
rect 1083 554 1129 566
rect 1241 742 1287 754
rect 1241 566 1247 742
rect 1281 566 1287 742
rect 1241 554 1287 566
rect 1399 742 1445 754
rect 1399 566 1405 742
rect 1439 566 1445 742
rect 1399 554 1445 566
rect 1557 742 1603 754
rect 1557 566 1563 742
rect 1597 566 1603 742
rect 1557 554 1603 566
rect 1715 742 1761 754
rect 1715 566 1721 742
rect 1755 566 1761 742
rect 1715 554 1761 566
rect 1873 742 1919 754
rect 1873 566 1879 742
rect 1913 566 1919 742
rect 1873 554 1919 566
rect 2031 742 2077 754
rect 2031 566 2037 742
rect 2071 566 2077 742
rect 2031 554 2077 566
rect 2189 742 2235 754
rect 2189 566 2195 742
rect 2229 566 2235 742
rect 2189 554 2235 566
rect -2179 507 -2087 513
rect -2179 473 -2167 507
rect -2099 473 -2087 507
rect -2179 467 -2087 473
rect -2021 507 -1929 513
rect -2021 473 -2009 507
rect -1941 473 -1929 507
rect -2021 467 -1929 473
rect -1863 507 -1771 513
rect -1863 473 -1851 507
rect -1783 473 -1771 507
rect -1863 467 -1771 473
rect -1705 507 -1613 513
rect -1705 473 -1693 507
rect -1625 473 -1613 507
rect -1705 467 -1613 473
rect -1547 507 -1455 513
rect -1547 473 -1535 507
rect -1467 473 -1455 507
rect -1547 467 -1455 473
rect -1389 507 -1297 513
rect -1389 473 -1377 507
rect -1309 473 -1297 507
rect -1389 467 -1297 473
rect -1231 507 -1139 513
rect -1231 473 -1219 507
rect -1151 473 -1139 507
rect -1231 467 -1139 473
rect -1073 507 -981 513
rect -1073 473 -1061 507
rect -993 473 -981 507
rect -1073 467 -981 473
rect -915 507 -823 513
rect -915 473 -903 507
rect -835 473 -823 507
rect -915 467 -823 473
rect -757 507 -665 513
rect -757 473 -745 507
rect -677 473 -665 507
rect -757 467 -665 473
rect -599 507 -507 513
rect -599 473 -587 507
rect -519 473 -507 507
rect -599 467 -507 473
rect -441 507 -349 513
rect -441 473 -429 507
rect -361 473 -349 507
rect -441 467 -349 473
rect -283 507 -191 513
rect -283 473 -271 507
rect -203 473 -191 507
rect -283 467 -191 473
rect -125 507 -33 513
rect -125 473 -113 507
rect -45 473 -33 507
rect -125 467 -33 473
rect 33 507 125 513
rect 33 473 45 507
rect 113 473 125 507
rect 33 467 125 473
rect 191 507 283 513
rect 191 473 203 507
rect 271 473 283 507
rect 191 467 283 473
rect 349 507 441 513
rect 349 473 361 507
rect 429 473 441 507
rect 349 467 441 473
rect 507 507 599 513
rect 507 473 519 507
rect 587 473 599 507
rect 507 467 599 473
rect 665 507 757 513
rect 665 473 677 507
rect 745 473 757 507
rect 665 467 757 473
rect 823 507 915 513
rect 823 473 835 507
rect 903 473 915 507
rect 823 467 915 473
rect 981 507 1073 513
rect 981 473 993 507
rect 1061 473 1073 507
rect 981 467 1073 473
rect 1139 507 1231 513
rect 1139 473 1151 507
rect 1219 473 1231 507
rect 1139 467 1231 473
rect 1297 507 1389 513
rect 1297 473 1309 507
rect 1377 473 1389 507
rect 1297 467 1389 473
rect 1455 507 1547 513
rect 1455 473 1467 507
rect 1535 473 1547 507
rect 1455 467 1547 473
rect 1613 507 1705 513
rect 1613 473 1625 507
rect 1693 473 1705 507
rect 1613 467 1705 473
rect 1771 507 1863 513
rect 1771 473 1783 507
rect 1851 473 1863 507
rect 1771 467 1863 473
rect 1929 507 2021 513
rect 1929 473 1941 507
rect 2009 473 2021 507
rect 1929 467 2021 473
rect 2087 507 2179 513
rect 2087 473 2099 507
rect 2167 473 2179 507
rect 2087 467 2179 473
rect -2179 399 -2087 405
rect -2179 365 -2167 399
rect -2099 365 -2087 399
rect -2179 359 -2087 365
rect -2021 399 -1929 405
rect -2021 365 -2009 399
rect -1941 365 -1929 399
rect -2021 359 -1929 365
rect -1863 399 -1771 405
rect -1863 365 -1851 399
rect -1783 365 -1771 399
rect -1863 359 -1771 365
rect -1705 399 -1613 405
rect -1705 365 -1693 399
rect -1625 365 -1613 399
rect -1705 359 -1613 365
rect -1547 399 -1455 405
rect -1547 365 -1535 399
rect -1467 365 -1455 399
rect -1547 359 -1455 365
rect -1389 399 -1297 405
rect -1389 365 -1377 399
rect -1309 365 -1297 399
rect -1389 359 -1297 365
rect -1231 399 -1139 405
rect -1231 365 -1219 399
rect -1151 365 -1139 399
rect -1231 359 -1139 365
rect -1073 399 -981 405
rect -1073 365 -1061 399
rect -993 365 -981 399
rect -1073 359 -981 365
rect -915 399 -823 405
rect -915 365 -903 399
rect -835 365 -823 399
rect -915 359 -823 365
rect -757 399 -665 405
rect -757 365 -745 399
rect -677 365 -665 399
rect -757 359 -665 365
rect -599 399 -507 405
rect -599 365 -587 399
rect -519 365 -507 399
rect -599 359 -507 365
rect -441 399 -349 405
rect -441 365 -429 399
rect -361 365 -349 399
rect -441 359 -349 365
rect -283 399 -191 405
rect -283 365 -271 399
rect -203 365 -191 399
rect -283 359 -191 365
rect -125 399 -33 405
rect -125 365 -113 399
rect -45 365 -33 399
rect -125 359 -33 365
rect 33 399 125 405
rect 33 365 45 399
rect 113 365 125 399
rect 33 359 125 365
rect 191 399 283 405
rect 191 365 203 399
rect 271 365 283 399
rect 191 359 283 365
rect 349 399 441 405
rect 349 365 361 399
rect 429 365 441 399
rect 349 359 441 365
rect 507 399 599 405
rect 507 365 519 399
rect 587 365 599 399
rect 507 359 599 365
rect 665 399 757 405
rect 665 365 677 399
rect 745 365 757 399
rect 665 359 757 365
rect 823 399 915 405
rect 823 365 835 399
rect 903 365 915 399
rect 823 359 915 365
rect 981 399 1073 405
rect 981 365 993 399
rect 1061 365 1073 399
rect 981 359 1073 365
rect 1139 399 1231 405
rect 1139 365 1151 399
rect 1219 365 1231 399
rect 1139 359 1231 365
rect 1297 399 1389 405
rect 1297 365 1309 399
rect 1377 365 1389 399
rect 1297 359 1389 365
rect 1455 399 1547 405
rect 1455 365 1467 399
rect 1535 365 1547 399
rect 1455 359 1547 365
rect 1613 399 1705 405
rect 1613 365 1625 399
rect 1693 365 1705 399
rect 1613 359 1705 365
rect 1771 399 1863 405
rect 1771 365 1783 399
rect 1851 365 1863 399
rect 1771 359 1863 365
rect 1929 399 2021 405
rect 1929 365 1941 399
rect 2009 365 2021 399
rect 1929 359 2021 365
rect 2087 399 2179 405
rect 2087 365 2099 399
rect 2167 365 2179 399
rect 2087 359 2179 365
rect -2235 306 -2189 318
rect -2235 130 -2229 306
rect -2195 130 -2189 306
rect -2235 118 -2189 130
rect -2077 306 -2031 318
rect -2077 130 -2071 306
rect -2037 130 -2031 306
rect -2077 118 -2031 130
rect -1919 306 -1873 318
rect -1919 130 -1913 306
rect -1879 130 -1873 306
rect -1919 118 -1873 130
rect -1761 306 -1715 318
rect -1761 130 -1755 306
rect -1721 130 -1715 306
rect -1761 118 -1715 130
rect -1603 306 -1557 318
rect -1603 130 -1597 306
rect -1563 130 -1557 306
rect -1603 118 -1557 130
rect -1445 306 -1399 318
rect -1445 130 -1439 306
rect -1405 130 -1399 306
rect -1445 118 -1399 130
rect -1287 306 -1241 318
rect -1287 130 -1281 306
rect -1247 130 -1241 306
rect -1287 118 -1241 130
rect -1129 306 -1083 318
rect -1129 130 -1123 306
rect -1089 130 -1083 306
rect -1129 118 -1083 130
rect -971 306 -925 318
rect -971 130 -965 306
rect -931 130 -925 306
rect -971 118 -925 130
rect -813 306 -767 318
rect -813 130 -807 306
rect -773 130 -767 306
rect -813 118 -767 130
rect -655 306 -609 318
rect -655 130 -649 306
rect -615 130 -609 306
rect -655 118 -609 130
rect -497 306 -451 318
rect -497 130 -491 306
rect -457 130 -451 306
rect -497 118 -451 130
rect -339 306 -293 318
rect -339 130 -333 306
rect -299 130 -293 306
rect -339 118 -293 130
rect -181 306 -135 318
rect -181 130 -175 306
rect -141 130 -135 306
rect -181 118 -135 130
rect -23 306 23 318
rect -23 130 -17 306
rect 17 130 23 306
rect -23 118 23 130
rect 135 306 181 318
rect 135 130 141 306
rect 175 130 181 306
rect 135 118 181 130
rect 293 306 339 318
rect 293 130 299 306
rect 333 130 339 306
rect 293 118 339 130
rect 451 306 497 318
rect 451 130 457 306
rect 491 130 497 306
rect 451 118 497 130
rect 609 306 655 318
rect 609 130 615 306
rect 649 130 655 306
rect 609 118 655 130
rect 767 306 813 318
rect 767 130 773 306
rect 807 130 813 306
rect 767 118 813 130
rect 925 306 971 318
rect 925 130 931 306
rect 965 130 971 306
rect 925 118 971 130
rect 1083 306 1129 318
rect 1083 130 1089 306
rect 1123 130 1129 306
rect 1083 118 1129 130
rect 1241 306 1287 318
rect 1241 130 1247 306
rect 1281 130 1287 306
rect 1241 118 1287 130
rect 1399 306 1445 318
rect 1399 130 1405 306
rect 1439 130 1445 306
rect 1399 118 1445 130
rect 1557 306 1603 318
rect 1557 130 1563 306
rect 1597 130 1603 306
rect 1557 118 1603 130
rect 1715 306 1761 318
rect 1715 130 1721 306
rect 1755 130 1761 306
rect 1715 118 1761 130
rect 1873 306 1919 318
rect 1873 130 1879 306
rect 1913 130 1919 306
rect 1873 118 1919 130
rect 2031 306 2077 318
rect 2031 130 2037 306
rect 2071 130 2077 306
rect 2031 118 2077 130
rect 2189 306 2235 318
rect 2189 130 2195 306
rect 2229 130 2235 306
rect 2189 118 2235 130
rect -2179 71 -2087 77
rect -2179 37 -2167 71
rect -2099 37 -2087 71
rect -2179 31 -2087 37
rect -2021 71 -1929 77
rect -2021 37 -2009 71
rect -1941 37 -1929 71
rect -2021 31 -1929 37
rect -1863 71 -1771 77
rect -1863 37 -1851 71
rect -1783 37 -1771 71
rect -1863 31 -1771 37
rect -1705 71 -1613 77
rect -1705 37 -1693 71
rect -1625 37 -1613 71
rect -1705 31 -1613 37
rect -1547 71 -1455 77
rect -1547 37 -1535 71
rect -1467 37 -1455 71
rect -1547 31 -1455 37
rect -1389 71 -1297 77
rect -1389 37 -1377 71
rect -1309 37 -1297 71
rect -1389 31 -1297 37
rect -1231 71 -1139 77
rect -1231 37 -1219 71
rect -1151 37 -1139 71
rect -1231 31 -1139 37
rect -1073 71 -981 77
rect -1073 37 -1061 71
rect -993 37 -981 71
rect -1073 31 -981 37
rect -915 71 -823 77
rect -915 37 -903 71
rect -835 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 835 71
rect 903 37 915 71
rect 823 31 915 37
rect 981 71 1073 77
rect 981 37 993 71
rect 1061 37 1073 71
rect 981 31 1073 37
rect 1139 71 1231 77
rect 1139 37 1151 71
rect 1219 37 1231 71
rect 1139 31 1231 37
rect 1297 71 1389 77
rect 1297 37 1309 71
rect 1377 37 1389 71
rect 1297 31 1389 37
rect 1455 71 1547 77
rect 1455 37 1467 71
rect 1535 37 1547 71
rect 1455 31 1547 37
rect 1613 71 1705 77
rect 1613 37 1625 71
rect 1693 37 1705 71
rect 1613 31 1705 37
rect 1771 71 1863 77
rect 1771 37 1783 71
rect 1851 37 1863 71
rect 1771 31 1863 37
rect 1929 71 2021 77
rect 1929 37 1941 71
rect 2009 37 2021 71
rect 1929 31 2021 37
rect 2087 71 2179 77
rect 2087 37 2099 71
rect 2167 37 2179 71
rect 2087 31 2179 37
rect -2179 -37 -2087 -31
rect -2179 -71 -2167 -37
rect -2099 -71 -2087 -37
rect -2179 -77 -2087 -71
rect -2021 -37 -1929 -31
rect -2021 -71 -2009 -37
rect -1941 -71 -1929 -37
rect -2021 -77 -1929 -71
rect -1863 -37 -1771 -31
rect -1863 -71 -1851 -37
rect -1783 -71 -1771 -37
rect -1863 -77 -1771 -71
rect -1705 -37 -1613 -31
rect -1705 -71 -1693 -37
rect -1625 -71 -1613 -37
rect -1705 -77 -1613 -71
rect -1547 -37 -1455 -31
rect -1547 -71 -1535 -37
rect -1467 -71 -1455 -37
rect -1547 -77 -1455 -71
rect -1389 -37 -1297 -31
rect -1389 -71 -1377 -37
rect -1309 -71 -1297 -37
rect -1389 -77 -1297 -71
rect -1231 -37 -1139 -31
rect -1231 -71 -1219 -37
rect -1151 -71 -1139 -37
rect -1231 -77 -1139 -71
rect -1073 -37 -981 -31
rect -1073 -71 -1061 -37
rect -993 -71 -981 -37
rect -1073 -77 -981 -71
rect -915 -37 -823 -31
rect -915 -71 -903 -37
rect -835 -71 -823 -37
rect -915 -77 -823 -71
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect 823 -37 915 -31
rect 823 -71 835 -37
rect 903 -71 915 -37
rect 823 -77 915 -71
rect 981 -37 1073 -31
rect 981 -71 993 -37
rect 1061 -71 1073 -37
rect 981 -77 1073 -71
rect 1139 -37 1231 -31
rect 1139 -71 1151 -37
rect 1219 -71 1231 -37
rect 1139 -77 1231 -71
rect 1297 -37 1389 -31
rect 1297 -71 1309 -37
rect 1377 -71 1389 -37
rect 1297 -77 1389 -71
rect 1455 -37 1547 -31
rect 1455 -71 1467 -37
rect 1535 -71 1547 -37
rect 1455 -77 1547 -71
rect 1613 -37 1705 -31
rect 1613 -71 1625 -37
rect 1693 -71 1705 -37
rect 1613 -77 1705 -71
rect 1771 -37 1863 -31
rect 1771 -71 1783 -37
rect 1851 -71 1863 -37
rect 1771 -77 1863 -71
rect 1929 -37 2021 -31
rect 1929 -71 1941 -37
rect 2009 -71 2021 -37
rect 1929 -77 2021 -71
rect 2087 -37 2179 -31
rect 2087 -71 2099 -37
rect 2167 -71 2179 -37
rect 2087 -77 2179 -71
rect -2235 -130 -2189 -118
rect -2235 -306 -2229 -130
rect -2195 -306 -2189 -130
rect -2235 -318 -2189 -306
rect -2077 -130 -2031 -118
rect -2077 -306 -2071 -130
rect -2037 -306 -2031 -130
rect -2077 -318 -2031 -306
rect -1919 -130 -1873 -118
rect -1919 -306 -1913 -130
rect -1879 -306 -1873 -130
rect -1919 -318 -1873 -306
rect -1761 -130 -1715 -118
rect -1761 -306 -1755 -130
rect -1721 -306 -1715 -130
rect -1761 -318 -1715 -306
rect -1603 -130 -1557 -118
rect -1603 -306 -1597 -130
rect -1563 -306 -1557 -130
rect -1603 -318 -1557 -306
rect -1445 -130 -1399 -118
rect -1445 -306 -1439 -130
rect -1405 -306 -1399 -130
rect -1445 -318 -1399 -306
rect -1287 -130 -1241 -118
rect -1287 -306 -1281 -130
rect -1247 -306 -1241 -130
rect -1287 -318 -1241 -306
rect -1129 -130 -1083 -118
rect -1129 -306 -1123 -130
rect -1089 -306 -1083 -130
rect -1129 -318 -1083 -306
rect -971 -130 -925 -118
rect -971 -306 -965 -130
rect -931 -306 -925 -130
rect -971 -318 -925 -306
rect -813 -130 -767 -118
rect -813 -306 -807 -130
rect -773 -306 -767 -130
rect -813 -318 -767 -306
rect -655 -130 -609 -118
rect -655 -306 -649 -130
rect -615 -306 -609 -130
rect -655 -318 -609 -306
rect -497 -130 -451 -118
rect -497 -306 -491 -130
rect -457 -306 -451 -130
rect -497 -318 -451 -306
rect -339 -130 -293 -118
rect -339 -306 -333 -130
rect -299 -306 -293 -130
rect -339 -318 -293 -306
rect -181 -130 -135 -118
rect -181 -306 -175 -130
rect -141 -306 -135 -130
rect -181 -318 -135 -306
rect -23 -130 23 -118
rect -23 -306 -17 -130
rect 17 -306 23 -130
rect -23 -318 23 -306
rect 135 -130 181 -118
rect 135 -306 141 -130
rect 175 -306 181 -130
rect 135 -318 181 -306
rect 293 -130 339 -118
rect 293 -306 299 -130
rect 333 -306 339 -130
rect 293 -318 339 -306
rect 451 -130 497 -118
rect 451 -306 457 -130
rect 491 -306 497 -130
rect 451 -318 497 -306
rect 609 -130 655 -118
rect 609 -306 615 -130
rect 649 -306 655 -130
rect 609 -318 655 -306
rect 767 -130 813 -118
rect 767 -306 773 -130
rect 807 -306 813 -130
rect 767 -318 813 -306
rect 925 -130 971 -118
rect 925 -306 931 -130
rect 965 -306 971 -130
rect 925 -318 971 -306
rect 1083 -130 1129 -118
rect 1083 -306 1089 -130
rect 1123 -306 1129 -130
rect 1083 -318 1129 -306
rect 1241 -130 1287 -118
rect 1241 -306 1247 -130
rect 1281 -306 1287 -130
rect 1241 -318 1287 -306
rect 1399 -130 1445 -118
rect 1399 -306 1405 -130
rect 1439 -306 1445 -130
rect 1399 -318 1445 -306
rect 1557 -130 1603 -118
rect 1557 -306 1563 -130
rect 1597 -306 1603 -130
rect 1557 -318 1603 -306
rect 1715 -130 1761 -118
rect 1715 -306 1721 -130
rect 1755 -306 1761 -130
rect 1715 -318 1761 -306
rect 1873 -130 1919 -118
rect 1873 -306 1879 -130
rect 1913 -306 1919 -130
rect 1873 -318 1919 -306
rect 2031 -130 2077 -118
rect 2031 -306 2037 -130
rect 2071 -306 2077 -130
rect 2031 -318 2077 -306
rect 2189 -130 2235 -118
rect 2189 -306 2195 -130
rect 2229 -306 2235 -130
rect 2189 -318 2235 -306
rect -2179 -365 -2087 -359
rect -2179 -399 -2167 -365
rect -2099 -399 -2087 -365
rect -2179 -405 -2087 -399
rect -2021 -365 -1929 -359
rect -2021 -399 -2009 -365
rect -1941 -399 -1929 -365
rect -2021 -405 -1929 -399
rect -1863 -365 -1771 -359
rect -1863 -399 -1851 -365
rect -1783 -399 -1771 -365
rect -1863 -405 -1771 -399
rect -1705 -365 -1613 -359
rect -1705 -399 -1693 -365
rect -1625 -399 -1613 -365
rect -1705 -405 -1613 -399
rect -1547 -365 -1455 -359
rect -1547 -399 -1535 -365
rect -1467 -399 -1455 -365
rect -1547 -405 -1455 -399
rect -1389 -365 -1297 -359
rect -1389 -399 -1377 -365
rect -1309 -399 -1297 -365
rect -1389 -405 -1297 -399
rect -1231 -365 -1139 -359
rect -1231 -399 -1219 -365
rect -1151 -399 -1139 -365
rect -1231 -405 -1139 -399
rect -1073 -365 -981 -359
rect -1073 -399 -1061 -365
rect -993 -399 -981 -365
rect -1073 -405 -981 -399
rect -915 -365 -823 -359
rect -915 -399 -903 -365
rect -835 -399 -823 -365
rect -915 -405 -823 -399
rect -757 -365 -665 -359
rect -757 -399 -745 -365
rect -677 -399 -665 -365
rect -757 -405 -665 -399
rect -599 -365 -507 -359
rect -599 -399 -587 -365
rect -519 -399 -507 -365
rect -599 -405 -507 -399
rect -441 -365 -349 -359
rect -441 -399 -429 -365
rect -361 -399 -349 -365
rect -441 -405 -349 -399
rect -283 -365 -191 -359
rect -283 -399 -271 -365
rect -203 -399 -191 -365
rect -283 -405 -191 -399
rect -125 -365 -33 -359
rect -125 -399 -113 -365
rect -45 -399 -33 -365
rect -125 -405 -33 -399
rect 33 -365 125 -359
rect 33 -399 45 -365
rect 113 -399 125 -365
rect 33 -405 125 -399
rect 191 -365 283 -359
rect 191 -399 203 -365
rect 271 -399 283 -365
rect 191 -405 283 -399
rect 349 -365 441 -359
rect 349 -399 361 -365
rect 429 -399 441 -365
rect 349 -405 441 -399
rect 507 -365 599 -359
rect 507 -399 519 -365
rect 587 -399 599 -365
rect 507 -405 599 -399
rect 665 -365 757 -359
rect 665 -399 677 -365
rect 745 -399 757 -365
rect 665 -405 757 -399
rect 823 -365 915 -359
rect 823 -399 835 -365
rect 903 -399 915 -365
rect 823 -405 915 -399
rect 981 -365 1073 -359
rect 981 -399 993 -365
rect 1061 -399 1073 -365
rect 981 -405 1073 -399
rect 1139 -365 1231 -359
rect 1139 -399 1151 -365
rect 1219 -399 1231 -365
rect 1139 -405 1231 -399
rect 1297 -365 1389 -359
rect 1297 -399 1309 -365
rect 1377 -399 1389 -365
rect 1297 -405 1389 -399
rect 1455 -365 1547 -359
rect 1455 -399 1467 -365
rect 1535 -399 1547 -365
rect 1455 -405 1547 -399
rect 1613 -365 1705 -359
rect 1613 -399 1625 -365
rect 1693 -399 1705 -365
rect 1613 -405 1705 -399
rect 1771 -365 1863 -359
rect 1771 -399 1783 -365
rect 1851 -399 1863 -365
rect 1771 -405 1863 -399
rect 1929 -365 2021 -359
rect 1929 -399 1941 -365
rect 2009 -399 2021 -365
rect 1929 -405 2021 -399
rect 2087 -365 2179 -359
rect 2087 -399 2099 -365
rect 2167 -399 2179 -365
rect 2087 -405 2179 -399
rect -2179 -473 -2087 -467
rect -2179 -507 -2167 -473
rect -2099 -507 -2087 -473
rect -2179 -513 -2087 -507
rect -2021 -473 -1929 -467
rect -2021 -507 -2009 -473
rect -1941 -507 -1929 -473
rect -2021 -513 -1929 -507
rect -1863 -473 -1771 -467
rect -1863 -507 -1851 -473
rect -1783 -507 -1771 -473
rect -1863 -513 -1771 -507
rect -1705 -473 -1613 -467
rect -1705 -507 -1693 -473
rect -1625 -507 -1613 -473
rect -1705 -513 -1613 -507
rect -1547 -473 -1455 -467
rect -1547 -507 -1535 -473
rect -1467 -507 -1455 -473
rect -1547 -513 -1455 -507
rect -1389 -473 -1297 -467
rect -1389 -507 -1377 -473
rect -1309 -507 -1297 -473
rect -1389 -513 -1297 -507
rect -1231 -473 -1139 -467
rect -1231 -507 -1219 -473
rect -1151 -507 -1139 -473
rect -1231 -513 -1139 -507
rect -1073 -473 -981 -467
rect -1073 -507 -1061 -473
rect -993 -507 -981 -473
rect -1073 -513 -981 -507
rect -915 -473 -823 -467
rect -915 -507 -903 -473
rect -835 -507 -823 -473
rect -915 -513 -823 -507
rect -757 -473 -665 -467
rect -757 -507 -745 -473
rect -677 -507 -665 -473
rect -757 -513 -665 -507
rect -599 -473 -507 -467
rect -599 -507 -587 -473
rect -519 -507 -507 -473
rect -599 -513 -507 -507
rect -441 -473 -349 -467
rect -441 -507 -429 -473
rect -361 -507 -349 -473
rect -441 -513 -349 -507
rect -283 -473 -191 -467
rect -283 -507 -271 -473
rect -203 -507 -191 -473
rect -283 -513 -191 -507
rect -125 -473 -33 -467
rect -125 -507 -113 -473
rect -45 -507 -33 -473
rect -125 -513 -33 -507
rect 33 -473 125 -467
rect 33 -507 45 -473
rect 113 -507 125 -473
rect 33 -513 125 -507
rect 191 -473 283 -467
rect 191 -507 203 -473
rect 271 -507 283 -473
rect 191 -513 283 -507
rect 349 -473 441 -467
rect 349 -507 361 -473
rect 429 -507 441 -473
rect 349 -513 441 -507
rect 507 -473 599 -467
rect 507 -507 519 -473
rect 587 -507 599 -473
rect 507 -513 599 -507
rect 665 -473 757 -467
rect 665 -507 677 -473
rect 745 -507 757 -473
rect 665 -513 757 -507
rect 823 -473 915 -467
rect 823 -507 835 -473
rect 903 -507 915 -473
rect 823 -513 915 -507
rect 981 -473 1073 -467
rect 981 -507 993 -473
rect 1061 -507 1073 -473
rect 981 -513 1073 -507
rect 1139 -473 1231 -467
rect 1139 -507 1151 -473
rect 1219 -507 1231 -473
rect 1139 -513 1231 -507
rect 1297 -473 1389 -467
rect 1297 -507 1309 -473
rect 1377 -507 1389 -473
rect 1297 -513 1389 -507
rect 1455 -473 1547 -467
rect 1455 -507 1467 -473
rect 1535 -507 1547 -473
rect 1455 -513 1547 -507
rect 1613 -473 1705 -467
rect 1613 -507 1625 -473
rect 1693 -507 1705 -473
rect 1613 -513 1705 -507
rect 1771 -473 1863 -467
rect 1771 -507 1783 -473
rect 1851 -507 1863 -473
rect 1771 -513 1863 -507
rect 1929 -473 2021 -467
rect 1929 -507 1941 -473
rect 2009 -507 2021 -473
rect 1929 -513 2021 -507
rect 2087 -473 2179 -467
rect 2087 -507 2099 -473
rect 2167 -507 2179 -473
rect 2087 -513 2179 -507
rect -2235 -566 -2189 -554
rect -2235 -742 -2229 -566
rect -2195 -742 -2189 -566
rect -2235 -754 -2189 -742
rect -2077 -566 -2031 -554
rect -2077 -742 -2071 -566
rect -2037 -742 -2031 -566
rect -2077 -754 -2031 -742
rect -1919 -566 -1873 -554
rect -1919 -742 -1913 -566
rect -1879 -742 -1873 -566
rect -1919 -754 -1873 -742
rect -1761 -566 -1715 -554
rect -1761 -742 -1755 -566
rect -1721 -742 -1715 -566
rect -1761 -754 -1715 -742
rect -1603 -566 -1557 -554
rect -1603 -742 -1597 -566
rect -1563 -742 -1557 -566
rect -1603 -754 -1557 -742
rect -1445 -566 -1399 -554
rect -1445 -742 -1439 -566
rect -1405 -742 -1399 -566
rect -1445 -754 -1399 -742
rect -1287 -566 -1241 -554
rect -1287 -742 -1281 -566
rect -1247 -742 -1241 -566
rect -1287 -754 -1241 -742
rect -1129 -566 -1083 -554
rect -1129 -742 -1123 -566
rect -1089 -742 -1083 -566
rect -1129 -754 -1083 -742
rect -971 -566 -925 -554
rect -971 -742 -965 -566
rect -931 -742 -925 -566
rect -971 -754 -925 -742
rect -813 -566 -767 -554
rect -813 -742 -807 -566
rect -773 -742 -767 -566
rect -813 -754 -767 -742
rect -655 -566 -609 -554
rect -655 -742 -649 -566
rect -615 -742 -609 -566
rect -655 -754 -609 -742
rect -497 -566 -451 -554
rect -497 -742 -491 -566
rect -457 -742 -451 -566
rect -497 -754 -451 -742
rect -339 -566 -293 -554
rect -339 -742 -333 -566
rect -299 -742 -293 -566
rect -339 -754 -293 -742
rect -181 -566 -135 -554
rect -181 -742 -175 -566
rect -141 -742 -135 -566
rect -181 -754 -135 -742
rect -23 -566 23 -554
rect -23 -742 -17 -566
rect 17 -742 23 -566
rect -23 -754 23 -742
rect 135 -566 181 -554
rect 135 -742 141 -566
rect 175 -742 181 -566
rect 135 -754 181 -742
rect 293 -566 339 -554
rect 293 -742 299 -566
rect 333 -742 339 -566
rect 293 -754 339 -742
rect 451 -566 497 -554
rect 451 -742 457 -566
rect 491 -742 497 -566
rect 451 -754 497 -742
rect 609 -566 655 -554
rect 609 -742 615 -566
rect 649 -742 655 -566
rect 609 -754 655 -742
rect 767 -566 813 -554
rect 767 -742 773 -566
rect 807 -742 813 -566
rect 767 -754 813 -742
rect 925 -566 971 -554
rect 925 -742 931 -566
rect 965 -742 971 -566
rect 925 -754 971 -742
rect 1083 -566 1129 -554
rect 1083 -742 1089 -566
rect 1123 -742 1129 -566
rect 1083 -754 1129 -742
rect 1241 -566 1287 -554
rect 1241 -742 1247 -566
rect 1281 -742 1287 -566
rect 1241 -754 1287 -742
rect 1399 -566 1445 -554
rect 1399 -742 1405 -566
rect 1439 -742 1445 -566
rect 1399 -754 1445 -742
rect 1557 -566 1603 -554
rect 1557 -742 1563 -566
rect 1597 -742 1603 -566
rect 1557 -754 1603 -742
rect 1715 -566 1761 -554
rect 1715 -742 1721 -566
rect 1755 -742 1761 -566
rect 1715 -754 1761 -742
rect 1873 -566 1919 -554
rect 1873 -742 1879 -566
rect 1913 -742 1919 -566
rect 1873 -754 1919 -742
rect 2031 -566 2077 -554
rect 2031 -742 2037 -566
rect 2071 -742 2077 -566
rect 2031 -754 2077 -742
rect 2189 -566 2235 -554
rect 2189 -742 2195 -566
rect 2229 -742 2235 -566
rect 2189 -754 2235 -742
rect -2179 -801 -2087 -795
rect -2179 -835 -2167 -801
rect -2099 -835 -2087 -801
rect -2179 -841 -2087 -835
rect -2021 -801 -1929 -795
rect -2021 -835 -2009 -801
rect -1941 -835 -1929 -801
rect -2021 -841 -1929 -835
rect -1863 -801 -1771 -795
rect -1863 -835 -1851 -801
rect -1783 -835 -1771 -801
rect -1863 -841 -1771 -835
rect -1705 -801 -1613 -795
rect -1705 -835 -1693 -801
rect -1625 -835 -1613 -801
rect -1705 -841 -1613 -835
rect -1547 -801 -1455 -795
rect -1547 -835 -1535 -801
rect -1467 -835 -1455 -801
rect -1547 -841 -1455 -835
rect -1389 -801 -1297 -795
rect -1389 -835 -1377 -801
rect -1309 -835 -1297 -801
rect -1389 -841 -1297 -835
rect -1231 -801 -1139 -795
rect -1231 -835 -1219 -801
rect -1151 -835 -1139 -801
rect -1231 -841 -1139 -835
rect -1073 -801 -981 -795
rect -1073 -835 -1061 -801
rect -993 -835 -981 -801
rect -1073 -841 -981 -835
rect -915 -801 -823 -795
rect -915 -835 -903 -801
rect -835 -835 -823 -801
rect -915 -841 -823 -835
rect -757 -801 -665 -795
rect -757 -835 -745 -801
rect -677 -835 -665 -801
rect -757 -841 -665 -835
rect -599 -801 -507 -795
rect -599 -835 -587 -801
rect -519 -835 -507 -801
rect -599 -841 -507 -835
rect -441 -801 -349 -795
rect -441 -835 -429 -801
rect -361 -835 -349 -801
rect -441 -841 -349 -835
rect -283 -801 -191 -795
rect -283 -835 -271 -801
rect -203 -835 -191 -801
rect -283 -841 -191 -835
rect -125 -801 -33 -795
rect -125 -835 -113 -801
rect -45 -835 -33 -801
rect -125 -841 -33 -835
rect 33 -801 125 -795
rect 33 -835 45 -801
rect 113 -835 125 -801
rect 33 -841 125 -835
rect 191 -801 283 -795
rect 191 -835 203 -801
rect 271 -835 283 -801
rect 191 -841 283 -835
rect 349 -801 441 -795
rect 349 -835 361 -801
rect 429 -835 441 -801
rect 349 -841 441 -835
rect 507 -801 599 -795
rect 507 -835 519 -801
rect 587 -835 599 -801
rect 507 -841 599 -835
rect 665 -801 757 -795
rect 665 -835 677 -801
rect 745 -835 757 -801
rect 665 -841 757 -835
rect 823 -801 915 -795
rect 823 -835 835 -801
rect 903 -835 915 -801
rect 823 -841 915 -835
rect 981 -801 1073 -795
rect 981 -835 993 -801
rect 1061 -835 1073 -801
rect 981 -841 1073 -835
rect 1139 -801 1231 -795
rect 1139 -835 1151 -801
rect 1219 -835 1231 -801
rect 1139 -841 1231 -835
rect 1297 -801 1389 -795
rect 1297 -835 1309 -801
rect 1377 -835 1389 -801
rect 1297 -841 1389 -835
rect 1455 -801 1547 -795
rect 1455 -835 1467 -801
rect 1535 -835 1547 -801
rect 1455 -841 1547 -835
rect 1613 -801 1705 -795
rect 1613 -835 1625 -801
rect 1693 -835 1705 -801
rect 1613 -841 1705 -835
rect 1771 -801 1863 -795
rect 1771 -835 1783 -801
rect 1851 -835 1863 -801
rect 1771 -841 1863 -835
rect 1929 -801 2021 -795
rect 1929 -835 1941 -801
rect 2009 -835 2021 -801
rect 1929 -841 2021 -835
rect 2087 -801 2179 -795
rect 2087 -835 2099 -801
rect 2167 -835 2179 -801
rect 2087 -841 2179 -835
rect -2179 -909 -2087 -903
rect -2179 -943 -2167 -909
rect -2099 -943 -2087 -909
rect -2179 -949 -2087 -943
rect -2021 -909 -1929 -903
rect -2021 -943 -2009 -909
rect -1941 -943 -1929 -909
rect -2021 -949 -1929 -943
rect -1863 -909 -1771 -903
rect -1863 -943 -1851 -909
rect -1783 -943 -1771 -909
rect -1863 -949 -1771 -943
rect -1705 -909 -1613 -903
rect -1705 -943 -1693 -909
rect -1625 -943 -1613 -909
rect -1705 -949 -1613 -943
rect -1547 -909 -1455 -903
rect -1547 -943 -1535 -909
rect -1467 -943 -1455 -909
rect -1547 -949 -1455 -943
rect -1389 -909 -1297 -903
rect -1389 -943 -1377 -909
rect -1309 -943 -1297 -909
rect -1389 -949 -1297 -943
rect -1231 -909 -1139 -903
rect -1231 -943 -1219 -909
rect -1151 -943 -1139 -909
rect -1231 -949 -1139 -943
rect -1073 -909 -981 -903
rect -1073 -943 -1061 -909
rect -993 -943 -981 -909
rect -1073 -949 -981 -943
rect -915 -909 -823 -903
rect -915 -943 -903 -909
rect -835 -943 -823 -909
rect -915 -949 -823 -943
rect -757 -909 -665 -903
rect -757 -943 -745 -909
rect -677 -943 -665 -909
rect -757 -949 -665 -943
rect -599 -909 -507 -903
rect -599 -943 -587 -909
rect -519 -943 -507 -909
rect -599 -949 -507 -943
rect -441 -909 -349 -903
rect -441 -943 -429 -909
rect -361 -943 -349 -909
rect -441 -949 -349 -943
rect -283 -909 -191 -903
rect -283 -943 -271 -909
rect -203 -943 -191 -909
rect -283 -949 -191 -943
rect -125 -909 -33 -903
rect -125 -943 -113 -909
rect -45 -943 -33 -909
rect -125 -949 -33 -943
rect 33 -909 125 -903
rect 33 -943 45 -909
rect 113 -943 125 -909
rect 33 -949 125 -943
rect 191 -909 283 -903
rect 191 -943 203 -909
rect 271 -943 283 -909
rect 191 -949 283 -943
rect 349 -909 441 -903
rect 349 -943 361 -909
rect 429 -943 441 -909
rect 349 -949 441 -943
rect 507 -909 599 -903
rect 507 -943 519 -909
rect 587 -943 599 -909
rect 507 -949 599 -943
rect 665 -909 757 -903
rect 665 -943 677 -909
rect 745 -943 757 -909
rect 665 -949 757 -943
rect 823 -909 915 -903
rect 823 -943 835 -909
rect 903 -943 915 -909
rect 823 -949 915 -943
rect 981 -909 1073 -903
rect 981 -943 993 -909
rect 1061 -943 1073 -909
rect 981 -949 1073 -943
rect 1139 -909 1231 -903
rect 1139 -943 1151 -909
rect 1219 -943 1231 -909
rect 1139 -949 1231 -943
rect 1297 -909 1389 -903
rect 1297 -943 1309 -909
rect 1377 -943 1389 -909
rect 1297 -949 1389 -943
rect 1455 -909 1547 -903
rect 1455 -943 1467 -909
rect 1535 -943 1547 -909
rect 1455 -949 1547 -943
rect 1613 -909 1705 -903
rect 1613 -943 1625 -909
rect 1693 -943 1705 -909
rect 1613 -949 1705 -943
rect 1771 -909 1863 -903
rect 1771 -943 1783 -909
rect 1851 -943 1863 -909
rect 1771 -949 1863 -943
rect 1929 -909 2021 -903
rect 1929 -943 1941 -909
rect 2009 -943 2021 -909
rect 1929 -949 2021 -943
rect 2087 -909 2179 -903
rect 2087 -943 2099 -909
rect 2167 -943 2179 -909
rect 2087 -949 2179 -943
rect -2235 -1002 -2189 -990
rect -2235 -1178 -2229 -1002
rect -2195 -1178 -2189 -1002
rect -2235 -1190 -2189 -1178
rect -2077 -1002 -2031 -990
rect -2077 -1178 -2071 -1002
rect -2037 -1178 -2031 -1002
rect -2077 -1190 -2031 -1178
rect -1919 -1002 -1873 -990
rect -1919 -1178 -1913 -1002
rect -1879 -1178 -1873 -1002
rect -1919 -1190 -1873 -1178
rect -1761 -1002 -1715 -990
rect -1761 -1178 -1755 -1002
rect -1721 -1178 -1715 -1002
rect -1761 -1190 -1715 -1178
rect -1603 -1002 -1557 -990
rect -1603 -1178 -1597 -1002
rect -1563 -1178 -1557 -1002
rect -1603 -1190 -1557 -1178
rect -1445 -1002 -1399 -990
rect -1445 -1178 -1439 -1002
rect -1405 -1178 -1399 -1002
rect -1445 -1190 -1399 -1178
rect -1287 -1002 -1241 -990
rect -1287 -1178 -1281 -1002
rect -1247 -1178 -1241 -1002
rect -1287 -1190 -1241 -1178
rect -1129 -1002 -1083 -990
rect -1129 -1178 -1123 -1002
rect -1089 -1178 -1083 -1002
rect -1129 -1190 -1083 -1178
rect -971 -1002 -925 -990
rect -971 -1178 -965 -1002
rect -931 -1178 -925 -1002
rect -971 -1190 -925 -1178
rect -813 -1002 -767 -990
rect -813 -1178 -807 -1002
rect -773 -1178 -767 -1002
rect -813 -1190 -767 -1178
rect -655 -1002 -609 -990
rect -655 -1178 -649 -1002
rect -615 -1178 -609 -1002
rect -655 -1190 -609 -1178
rect -497 -1002 -451 -990
rect -497 -1178 -491 -1002
rect -457 -1178 -451 -1002
rect -497 -1190 -451 -1178
rect -339 -1002 -293 -990
rect -339 -1178 -333 -1002
rect -299 -1178 -293 -1002
rect -339 -1190 -293 -1178
rect -181 -1002 -135 -990
rect -181 -1178 -175 -1002
rect -141 -1178 -135 -1002
rect -181 -1190 -135 -1178
rect -23 -1002 23 -990
rect -23 -1178 -17 -1002
rect 17 -1178 23 -1002
rect -23 -1190 23 -1178
rect 135 -1002 181 -990
rect 135 -1178 141 -1002
rect 175 -1178 181 -1002
rect 135 -1190 181 -1178
rect 293 -1002 339 -990
rect 293 -1178 299 -1002
rect 333 -1178 339 -1002
rect 293 -1190 339 -1178
rect 451 -1002 497 -990
rect 451 -1178 457 -1002
rect 491 -1178 497 -1002
rect 451 -1190 497 -1178
rect 609 -1002 655 -990
rect 609 -1178 615 -1002
rect 649 -1178 655 -1002
rect 609 -1190 655 -1178
rect 767 -1002 813 -990
rect 767 -1178 773 -1002
rect 807 -1178 813 -1002
rect 767 -1190 813 -1178
rect 925 -1002 971 -990
rect 925 -1178 931 -1002
rect 965 -1178 971 -1002
rect 925 -1190 971 -1178
rect 1083 -1002 1129 -990
rect 1083 -1178 1089 -1002
rect 1123 -1178 1129 -1002
rect 1083 -1190 1129 -1178
rect 1241 -1002 1287 -990
rect 1241 -1178 1247 -1002
rect 1281 -1178 1287 -1002
rect 1241 -1190 1287 -1178
rect 1399 -1002 1445 -990
rect 1399 -1178 1405 -1002
rect 1439 -1178 1445 -1002
rect 1399 -1190 1445 -1178
rect 1557 -1002 1603 -990
rect 1557 -1178 1563 -1002
rect 1597 -1178 1603 -1002
rect 1557 -1190 1603 -1178
rect 1715 -1002 1761 -990
rect 1715 -1178 1721 -1002
rect 1755 -1178 1761 -1002
rect 1715 -1190 1761 -1178
rect 1873 -1002 1919 -990
rect 1873 -1178 1879 -1002
rect 1913 -1178 1919 -1002
rect 1873 -1190 1919 -1178
rect 2031 -1002 2077 -990
rect 2031 -1178 2037 -1002
rect 2071 -1178 2077 -1002
rect 2031 -1190 2077 -1178
rect 2189 -1002 2235 -990
rect 2189 -1178 2195 -1002
rect 2229 -1178 2235 -1002
rect 2189 -1190 2235 -1178
rect -2179 -1237 -2087 -1231
rect -2179 -1271 -2167 -1237
rect -2099 -1271 -2087 -1237
rect -2179 -1277 -2087 -1271
rect -2021 -1237 -1929 -1231
rect -2021 -1271 -2009 -1237
rect -1941 -1271 -1929 -1237
rect -2021 -1277 -1929 -1271
rect -1863 -1237 -1771 -1231
rect -1863 -1271 -1851 -1237
rect -1783 -1271 -1771 -1237
rect -1863 -1277 -1771 -1271
rect -1705 -1237 -1613 -1231
rect -1705 -1271 -1693 -1237
rect -1625 -1271 -1613 -1237
rect -1705 -1277 -1613 -1271
rect -1547 -1237 -1455 -1231
rect -1547 -1271 -1535 -1237
rect -1467 -1271 -1455 -1237
rect -1547 -1277 -1455 -1271
rect -1389 -1237 -1297 -1231
rect -1389 -1271 -1377 -1237
rect -1309 -1271 -1297 -1237
rect -1389 -1277 -1297 -1271
rect -1231 -1237 -1139 -1231
rect -1231 -1271 -1219 -1237
rect -1151 -1271 -1139 -1237
rect -1231 -1277 -1139 -1271
rect -1073 -1237 -981 -1231
rect -1073 -1271 -1061 -1237
rect -993 -1271 -981 -1237
rect -1073 -1277 -981 -1271
rect -915 -1237 -823 -1231
rect -915 -1271 -903 -1237
rect -835 -1271 -823 -1237
rect -915 -1277 -823 -1271
rect -757 -1237 -665 -1231
rect -757 -1271 -745 -1237
rect -677 -1271 -665 -1237
rect -757 -1277 -665 -1271
rect -599 -1237 -507 -1231
rect -599 -1271 -587 -1237
rect -519 -1271 -507 -1237
rect -599 -1277 -507 -1271
rect -441 -1237 -349 -1231
rect -441 -1271 -429 -1237
rect -361 -1271 -349 -1237
rect -441 -1277 -349 -1271
rect -283 -1237 -191 -1231
rect -283 -1271 -271 -1237
rect -203 -1271 -191 -1237
rect -283 -1277 -191 -1271
rect -125 -1237 -33 -1231
rect -125 -1271 -113 -1237
rect -45 -1271 -33 -1237
rect -125 -1277 -33 -1271
rect 33 -1237 125 -1231
rect 33 -1271 45 -1237
rect 113 -1271 125 -1237
rect 33 -1277 125 -1271
rect 191 -1237 283 -1231
rect 191 -1271 203 -1237
rect 271 -1271 283 -1237
rect 191 -1277 283 -1271
rect 349 -1237 441 -1231
rect 349 -1271 361 -1237
rect 429 -1271 441 -1237
rect 349 -1277 441 -1271
rect 507 -1237 599 -1231
rect 507 -1271 519 -1237
rect 587 -1271 599 -1237
rect 507 -1277 599 -1271
rect 665 -1237 757 -1231
rect 665 -1271 677 -1237
rect 745 -1271 757 -1237
rect 665 -1277 757 -1271
rect 823 -1237 915 -1231
rect 823 -1271 835 -1237
rect 903 -1271 915 -1237
rect 823 -1277 915 -1271
rect 981 -1237 1073 -1231
rect 981 -1271 993 -1237
rect 1061 -1271 1073 -1237
rect 981 -1277 1073 -1271
rect 1139 -1237 1231 -1231
rect 1139 -1271 1151 -1237
rect 1219 -1271 1231 -1237
rect 1139 -1277 1231 -1271
rect 1297 -1237 1389 -1231
rect 1297 -1271 1309 -1237
rect 1377 -1271 1389 -1237
rect 1297 -1277 1389 -1271
rect 1455 -1237 1547 -1231
rect 1455 -1271 1467 -1237
rect 1535 -1271 1547 -1237
rect 1455 -1277 1547 -1271
rect 1613 -1237 1705 -1231
rect 1613 -1271 1625 -1237
rect 1693 -1271 1705 -1237
rect 1613 -1277 1705 -1271
rect 1771 -1237 1863 -1231
rect 1771 -1271 1783 -1237
rect 1851 -1271 1863 -1237
rect 1771 -1277 1863 -1271
rect 1929 -1237 2021 -1231
rect 1929 -1271 1941 -1237
rect 2009 -1271 2021 -1237
rect 1929 -1277 2021 -1271
rect 2087 -1237 2179 -1231
rect 2087 -1271 2099 -1237
rect 2167 -1271 2179 -1237
rect 2087 -1277 2179 -1271
rect -2179 -1345 -2087 -1339
rect -2179 -1379 -2167 -1345
rect -2099 -1379 -2087 -1345
rect -2179 -1385 -2087 -1379
rect -2021 -1345 -1929 -1339
rect -2021 -1379 -2009 -1345
rect -1941 -1379 -1929 -1345
rect -2021 -1385 -1929 -1379
rect -1863 -1345 -1771 -1339
rect -1863 -1379 -1851 -1345
rect -1783 -1379 -1771 -1345
rect -1863 -1385 -1771 -1379
rect -1705 -1345 -1613 -1339
rect -1705 -1379 -1693 -1345
rect -1625 -1379 -1613 -1345
rect -1705 -1385 -1613 -1379
rect -1547 -1345 -1455 -1339
rect -1547 -1379 -1535 -1345
rect -1467 -1379 -1455 -1345
rect -1547 -1385 -1455 -1379
rect -1389 -1345 -1297 -1339
rect -1389 -1379 -1377 -1345
rect -1309 -1379 -1297 -1345
rect -1389 -1385 -1297 -1379
rect -1231 -1345 -1139 -1339
rect -1231 -1379 -1219 -1345
rect -1151 -1379 -1139 -1345
rect -1231 -1385 -1139 -1379
rect -1073 -1345 -981 -1339
rect -1073 -1379 -1061 -1345
rect -993 -1379 -981 -1345
rect -1073 -1385 -981 -1379
rect -915 -1345 -823 -1339
rect -915 -1379 -903 -1345
rect -835 -1379 -823 -1345
rect -915 -1385 -823 -1379
rect -757 -1345 -665 -1339
rect -757 -1379 -745 -1345
rect -677 -1379 -665 -1345
rect -757 -1385 -665 -1379
rect -599 -1345 -507 -1339
rect -599 -1379 -587 -1345
rect -519 -1379 -507 -1345
rect -599 -1385 -507 -1379
rect -441 -1345 -349 -1339
rect -441 -1379 -429 -1345
rect -361 -1379 -349 -1345
rect -441 -1385 -349 -1379
rect -283 -1345 -191 -1339
rect -283 -1379 -271 -1345
rect -203 -1379 -191 -1345
rect -283 -1385 -191 -1379
rect -125 -1345 -33 -1339
rect -125 -1379 -113 -1345
rect -45 -1379 -33 -1345
rect -125 -1385 -33 -1379
rect 33 -1345 125 -1339
rect 33 -1379 45 -1345
rect 113 -1379 125 -1345
rect 33 -1385 125 -1379
rect 191 -1345 283 -1339
rect 191 -1379 203 -1345
rect 271 -1379 283 -1345
rect 191 -1385 283 -1379
rect 349 -1345 441 -1339
rect 349 -1379 361 -1345
rect 429 -1379 441 -1345
rect 349 -1385 441 -1379
rect 507 -1345 599 -1339
rect 507 -1379 519 -1345
rect 587 -1379 599 -1345
rect 507 -1385 599 -1379
rect 665 -1345 757 -1339
rect 665 -1379 677 -1345
rect 745 -1379 757 -1345
rect 665 -1385 757 -1379
rect 823 -1345 915 -1339
rect 823 -1379 835 -1345
rect 903 -1379 915 -1345
rect 823 -1385 915 -1379
rect 981 -1345 1073 -1339
rect 981 -1379 993 -1345
rect 1061 -1379 1073 -1345
rect 981 -1385 1073 -1379
rect 1139 -1345 1231 -1339
rect 1139 -1379 1151 -1345
rect 1219 -1379 1231 -1345
rect 1139 -1385 1231 -1379
rect 1297 -1345 1389 -1339
rect 1297 -1379 1309 -1345
rect 1377 -1379 1389 -1345
rect 1297 -1385 1389 -1379
rect 1455 -1345 1547 -1339
rect 1455 -1379 1467 -1345
rect 1535 -1379 1547 -1345
rect 1455 -1385 1547 -1379
rect 1613 -1345 1705 -1339
rect 1613 -1379 1625 -1345
rect 1693 -1379 1705 -1345
rect 1613 -1385 1705 -1379
rect 1771 -1345 1863 -1339
rect 1771 -1379 1783 -1345
rect 1851 -1379 1863 -1345
rect 1771 -1385 1863 -1379
rect 1929 -1345 2021 -1339
rect 1929 -1379 1941 -1345
rect 2009 -1379 2021 -1345
rect 1929 -1385 2021 -1379
rect 2087 -1345 2179 -1339
rect 2087 -1379 2099 -1345
rect 2167 -1379 2179 -1345
rect 2087 -1385 2179 -1379
rect -2235 -1438 -2189 -1426
rect -2235 -1614 -2229 -1438
rect -2195 -1614 -2189 -1438
rect -2235 -1626 -2189 -1614
rect -2077 -1438 -2031 -1426
rect -2077 -1614 -2071 -1438
rect -2037 -1614 -2031 -1438
rect -2077 -1626 -2031 -1614
rect -1919 -1438 -1873 -1426
rect -1919 -1614 -1913 -1438
rect -1879 -1614 -1873 -1438
rect -1919 -1626 -1873 -1614
rect -1761 -1438 -1715 -1426
rect -1761 -1614 -1755 -1438
rect -1721 -1614 -1715 -1438
rect -1761 -1626 -1715 -1614
rect -1603 -1438 -1557 -1426
rect -1603 -1614 -1597 -1438
rect -1563 -1614 -1557 -1438
rect -1603 -1626 -1557 -1614
rect -1445 -1438 -1399 -1426
rect -1445 -1614 -1439 -1438
rect -1405 -1614 -1399 -1438
rect -1445 -1626 -1399 -1614
rect -1287 -1438 -1241 -1426
rect -1287 -1614 -1281 -1438
rect -1247 -1614 -1241 -1438
rect -1287 -1626 -1241 -1614
rect -1129 -1438 -1083 -1426
rect -1129 -1614 -1123 -1438
rect -1089 -1614 -1083 -1438
rect -1129 -1626 -1083 -1614
rect -971 -1438 -925 -1426
rect -971 -1614 -965 -1438
rect -931 -1614 -925 -1438
rect -971 -1626 -925 -1614
rect -813 -1438 -767 -1426
rect -813 -1614 -807 -1438
rect -773 -1614 -767 -1438
rect -813 -1626 -767 -1614
rect -655 -1438 -609 -1426
rect -655 -1614 -649 -1438
rect -615 -1614 -609 -1438
rect -655 -1626 -609 -1614
rect -497 -1438 -451 -1426
rect -497 -1614 -491 -1438
rect -457 -1614 -451 -1438
rect -497 -1626 -451 -1614
rect -339 -1438 -293 -1426
rect -339 -1614 -333 -1438
rect -299 -1614 -293 -1438
rect -339 -1626 -293 -1614
rect -181 -1438 -135 -1426
rect -181 -1614 -175 -1438
rect -141 -1614 -135 -1438
rect -181 -1626 -135 -1614
rect -23 -1438 23 -1426
rect -23 -1614 -17 -1438
rect 17 -1614 23 -1438
rect -23 -1626 23 -1614
rect 135 -1438 181 -1426
rect 135 -1614 141 -1438
rect 175 -1614 181 -1438
rect 135 -1626 181 -1614
rect 293 -1438 339 -1426
rect 293 -1614 299 -1438
rect 333 -1614 339 -1438
rect 293 -1626 339 -1614
rect 451 -1438 497 -1426
rect 451 -1614 457 -1438
rect 491 -1614 497 -1438
rect 451 -1626 497 -1614
rect 609 -1438 655 -1426
rect 609 -1614 615 -1438
rect 649 -1614 655 -1438
rect 609 -1626 655 -1614
rect 767 -1438 813 -1426
rect 767 -1614 773 -1438
rect 807 -1614 813 -1438
rect 767 -1626 813 -1614
rect 925 -1438 971 -1426
rect 925 -1614 931 -1438
rect 965 -1614 971 -1438
rect 925 -1626 971 -1614
rect 1083 -1438 1129 -1426
rect 1083 -1614 1089 -1438
rect 1123 -1614 1129 -1438
rect 1083 -1626 1129 -1614
rect 1241 -1438 1287 -1426
rect 1241 -1614 1247 -1438
rect 1281 -1614 1287 -1438
rect 1241 -1626 1287 -1614
rect 1399 -1438 1445 -1426
rect 1399 -1614 1405 -1438
rect 1439 -1614 1445 -1438
rect 1399 -1626 1445 -1614
rect 1557 -1438 1603 -1426
rect 1557 -1614 1563 -1438
rect 1597 -1614 1603 -1438
rect 1557 -1626 1603 -1614
rect 1715 -1438 1761 -1426
rect 1715 -1614 1721 -1438
rect 1755 -1614 1761 -1438
rect 1715 -1626 1761 -1614
rect 1873 -1438 1919 -1426
rect 1873 -1614 1879 -1438
rect 1913 -1614 1919 -1438
rect 1873 -1626 1919 -1614
rect 2031 -1438 2077 -1426
rect 2031 -1614 2037 -1438
rect 2071 -1614 2077 -1438
rect 2031 -1626 2077 -1614
rect 2189 -1438 2235 -1426
rect 2189 -1614 2195 -1438
rect 2229 -1614 2235 -1438
rect 2189 -1626 2235 -1614
rect -2179 -1673 -2087 -1667
rect -2179 -1707 -2167 -1673
rect -2099 -1707 -2087 -1673
rect -2179 -1713 -2087 -1707
rect -2021 -1673 -1929 -1667
rect -2021 -1707 -2009 -1673
rect -1941 -1707 -1929 -1673
rect -2021 -1713 -1929 -1707
rect -1863 -1673 -1771 -1667
rect -1863 -1707 -1851 -1673
rect -1783 -1707 -1771 -1673
rect -1863 -1713 -1771 -1707
rect -1705 -1673 -1613 -1667
rect -1705 -1707 -1693 -1673
rect -1625 -1707 -1613 -1673
rect -1705 -1713 -1613 -1707
rect -1547 -1673 -1455 -1667
rect -1547 -1707 -1535 -1673
rect -1467 -1707 -1455 -1673
rect -1547 -1713 -1455 -1707
rect -1389 -1673 -1297 -1667
rect -1389 -1707 -1377 -1673
rect -1309 -1707 -1297 -1673
rect -1389 -1713 -1297 -1707
rect -1231 -1673 -1139 -1667
rect -1231 -1707 -1219 -1673
rect -1151 -1707 -1139 -1673
rect -1231 -1713 -1139 -1707
rect -1073 -1673 -981 -1667
rect -1073 -1707 -1061 -1673
rect -993 -1707 -981 -1673
rect -1073 -1713 -981 -1707
rect -915 -1673 -823 -1667
rect -915 -1707 -903 -1673
rect -835 -1707 -823 -1673
rect -915 -1713 -823 -1707
rect -757 -1673 -665 -1667
rect -757 -1707 -745 -1673
rect -677 -1707 -665 -1673
rect -757 -1713 -665 -1707
rect -599 -1673 -507 -1667
rect -599 -1707 -587 -1673
rect -519 -1707 -507 -1673
rect -599 -1713 -507 -1707
rect -441 -1673 -349 -1667
rect -441 -1707 -429 -1673
rect -361 -1707 -349 -1673
rect -441 -1713 -349 -1707
rect -283 -1673 -191 -1667
rect -283 -1707 -271 -1673
rect -203 -1707 -191 -1673
rect -283 -1713 -191 -1707
rect -125 -1673 -33 -1667
rect -125 -1707 -113 -1673
rect -45 -1707 -33 -1673
rect -125 -1713 -33 -1707
rect 33 -1673 125 -1667
rect 33 -1707 45 -1673
rect 113 -1707 125 -1673
rect 33 -1713 125 -1707
rect 191 -1673 283 -1667
rect 191 -1707 203 -1673
rect 271 -1707 283 -1673
rect 191 -1713 283 -1707
rect 349 -1673 441 -1667
rect 349 -1707 361 -1673
rect 429 -1707 441 -1673
rect 349 -1713 441 -1707
rect 507 -1673 599 -1667
rect 507 -1707 519 -1673
rect 587 -1707 599 -1673
rect 507 -1713 599 -1707
rect 665 -1673 757 -1667
rect 665 -1707 677 -1673
rect 745 -1707 757 -1673
rect 665 -1713 757 -1707
rect 823 -1673 915 -1667
rect 823 -1707 835 -1673
rect 903 -1707 915 -1673
rect 823 -1713 915 -1707
rect 981 -1673 1073 -1667
rect 981 -1707 993 -1673
rect 1061 -1707 1073 -1673
rect 981 -1713 1073 -1707
rect 1139 -1673 1231 -1667
rect 1139 -1707 1151 -1673
rect 1219 -1707 1231 -1673
rect 1139 -1713 1231 -1707
rect 1297 -1673 1389 -1667
rect 1297 -1707 1309 -1673
rect 1377 -1707 1389 -1673
rect 1297 -1713 1389 -1707
rect 1455 -1673 1547 -1667
rect 1455 -1707 1467 -1673
rect 1535 -1707 1547 -1673
rect 1455 -1713 1547 -1707
rect 1613 -1673 1705 -1667
rect 1613 -1707 1625 -1673
rect 1693 -1707 1705 -1673
rect 1613 -1713 1705 -1707
rect 1771 -1673 1863 -1667
rect 1771 -1707 1783 -1673
rect 1851 -1707 1863 -1673
rect 1771 -1713 1863 -1707
rect 1929 -1673 2021 -1667
rect 1929 -1707 1941 -1673
rect 2009 -1707 2021 -1673
rect 1929 -1713 2021 -1707
rect 2087 -1673 2179 -1667
rect 2087 -1707 2099 -1673
rect 2167 -1707 2179 -1673
rect 2087 -1713 2179 -1707
rect -2179 -1781 -2087 -1775
rect -2179 -1815 -2167 -1781
rect -2099 -1815 -2087 -1781
rect -2179 -1821 -2087 -1815
rect -2021 -1781 -1929 -1775
rect -2021 -1815 -2009 -1781
rect -1941 -1815 -1929 -1781
rect -2021 -1821 -1929 -1815
rect -1863 -1781 -1771 -1775
rect -1863 -1815 -1851 -1781
rect -1783 -1815 -1771 -1781
rect -1863 -1821 -1771 -1815
rect -1705 -1781 -1613 -1775
rect -1705 -1815 -1693 -1781
rect -1625 -1815 -1613 -1781
rect -1705 -1821 -1613 -1815
rect -1547 -1781 -1455 -1775
rect -1547 -1815 -1535 -1781
rect -1467 -1815 -1455 -1781
rect -1547 -1821 -1455 -1815
rect -1389 -1781 -1297 -1775
rect -1389 -1815 -1377 -1781
rect -1309 -1815 -1297 -1781
rect -1389 -1821 -1297 -1815
rect -1231 -1781 -1139 -1775
rect -1231 -1815 -1219 -1781
rect -1151 -1815 -1139 -1781
rect -1231 -1821 -1139 -1815
rect -1073 -1781 -981 -1775
rect -1073 -1815 -1061 -1781
rect -993 -1815 -981 -1781
rect -1073 -1821 -981 -1815
rect -915 -1781 -823 -1775
rect -915 -1815 -903 -1781
rect -835 -1815 -823 -1781
rect -915 -1821 -823 -1815
rect -757 -1781 -665 -1775
rect -757 -1815 -745 -1781
rect -677 -1815 -665 -1781
rect -757 -1821 -665 -1815
rect -599 -1781 -507 -1775
rect -599 -1815 -587 -1781
rect -519 -1815 -507 -1781
rect -599 -1821 -507 -1815
rect -441 -1781 -349 -1775
rect -441 -1815 -429 -1781
rect -361 -1815 -349 -1781
rect -441 -1821 -349 -1815
rect -283 -1781 -191 -1775
rect -283 -1815 -271 -1781
rect -203 -1815 -191 -1781
rect -283 -1821 -191 -1815
rect -125 -1781 -33 -1775
rect -125 -1815 -113 -1781
rect -45 -1815 -33 -1781
rect -125 -1821 -33 -1815
rect 33 -1781 125 -1775
rect 33 -1815 45 -1781
rect 113 -1815 125 -1781
rect 33 -1821 125 -1815
rect 191 -1781 283 -1775
rect 191 -1815 203 -1781
rect 271 -1815 283 -1781
rect 191 -1821 283 -1815
rect 349 -1781 441 -1775
rect 349 -1815 361 -1781
rect 429 -1815 441 -1781
rect 349 -1821 441 -1815
rect 507 -1781 599 -1775
rect 507 -1815 519 -1781
rect 587 -1815 599 -1781
rect 507 -1821 599 -1815
rect 665 -1781 757 -1775
rect 665 -1815 677 -1781
rect 745 -1815 757 -1781
rect 665 -1821 757 -1815
rect 823 -1781 915 -1775
rect 823 -1815 835 -1781
rect 903 -1815 915 -1781
rect 823 -1821 915 -1815
rect 981 -1781 1073 -1775
rect 981 -1815 993 -1781
rect 1061 -1815 1073 -1781
rect 981 -1821 1073 -1815
rect 1139 -1781 1231 -1775
rect 1139 -1815 1151 -1781
rect 1219 -1815 1231 -1781
rect 1139 -1821 1231 -1815
rect 1297 -1781 1389 -1775
rect 1297 -1815 1309 -1781
rect 1377 -1815 1389 -1781
rect 1297 -1821 1389 -1815
rect 1455 -1781 1547 -1775
rect 1455 -1815 1467 -1781
rect 1535 -1815 1547 -1781
rect 1455 -1821 1547 -1815
rect 1613 -1781 1705 -1775
rect 1613 -1815 1625 -1781
rect 1693 -1815 1705 -1781
rect 1613 -1821 1705 -1815
rect 1771 -1781 1863 -1775
rect 1771 -1815 1783 -1781
rect 1851 -1815 1863 -1781
rect 1771 -1821 1863 -1815
rect 1929 -1781 2021 -1775
rect 1929 -1815 1941 -1781
rect 2009 -1815 2021 -1781
rect 1929 -1821 2021 -1815
rect 2087 -1781 2179 -1775
rect 2087 -1815 2099 -1781
rect 2167 -1815 2179 -1781
rect 2087 -1821 2179 -1815
rect -2235 -1874 -2189 -1862
rect -2235 -2050 -2229 -1874
rect -2195 -2050 -2189 -1874
rect -2235 -2062 -2189 -2050
rect -2077 -1874 -2031 -1862
rect -2077 -2050 -2071 -1874
rect -2037 -2050 -2031 -1874
rect -2077 -2062 -2031 -2050
rect -1919 -1874 -1873 -1862
rect -1919 -2050 -1913 -1874
rect -1879 -2050 -1873 -1874
rect -1919 -2062 -1873 -2050
rect -1761 -1874 -1715 -1862
rect -1761 -2050 -1755 -1874
rect -1721 -2050 -1715 -1874
rect -1761 -2062 -1715 -2050
rect -1603 -1874 -1557 -1862
rect -1603 -2050 -1597 -1874
rect -1563 -2050 -1557 -1874
rect -1603 -2062 -1557 -2050
rect -1445 -1874 -1399 -1862
rect -1445 -2050 -1439 -1874
rect -1405 -2050 -1399 -1874
rect -1445 -2062 -1399 -2050
rect -1287 -1874 -1241 -1862
rect -1287 -2050 -1281 -1874
rect -1247 -2050 -1241 -1874
rect -1287 -2062 -1241 -2050
rect -1129 -1874 -1083 -1862
rect -1129 -2050 -1123 -1874
rect -1089 -2050 -1083 -1874
rect -1129 -2062 -1083 -2050
rect -971 -1874 -925 -1862
rect -971 -2050 -965 -1874
rect -931 -2050 -925 -1874
rect -971 -2062 -925 -2050
rect -813 -1874 -767 -1862
rect -813 -2050 -807 -1874
rect -773 -2050 -767 -1874
rect -813 -2062 -767 -2050
rect -655 -1874 -609 -1862
rect -655 -2050 -649 -1874
rect -615 -2050 -609 -1874
rect -655 -2062 -609 -2050
rect -497 -1874 -451 -1862
rect -497 -2050 -491 -1874
rect -457 -2050 -451 -1874
rect -497 -2062 -451 -2050
rect -339 -1874 -293 -1862
rect -339 -2050 -333 -1874
rect -299 -2050 -293 -1874
rect -339 -2062 -293 -2050
rect -181 -1874 -135 -1862
rect -181 -2050 -175 -1874
rect -141 -2050 -135 -1874
rect -181 -2062 -135 -2050
rect -23 -1874 23 -1862
rect -23 -2050 -17 -1874
rect 17 -2050 23 -1874
rect -23 -2062 23 -2050
rect 135 -1874 181 -1862
rect 135 -2050 141 -1874
rect 175 -2050 181 -1874
rect 135 -2062 181 -2050
rect 293 -1874 339 -1862
rect 293 -2050 299 -1874
rect 333 -2050 339 -1874
rect 293 -2062 339 -2050
rect 451 -1874 497 -1862
rect 451 -2050 457 -1874
rect 491 -2050 497 -1874
rect 451 -2062 497 -2050
rect 609 -1874 655 -1862
rect 609 -2050 615 -1874
rect 649 -2050 655 -1874
rect 609 -2062 655 -2050
rect 767 -1874 813 -1862
rect 767 -2050 773 -1874
rect 807 -2050 813 -1874
rect 767 -2062 813 -2050
rect 925 -1874 971 -1862
rect 925 -2050 931 -1874
rect 965 -2050 971 -1874
rect 925 -2062 971 -2050
rect 1083 -1874 1129 -1862
rect 1083 -2050 1089 -1874
rect 1123 -2050 1129 -1874
rect 1083 -2062 1129 -2050
rect 1241 -1874 1287 -1862
rect 1241 -2050 1247 -1874
rect 1281 -2050 1287 -1874
rect 1241 -2062 1287 -2050
rect 1399 -1874 1445 -1862
rect 1399 -2050 1405 -1874
rect 1439 -2050 1445 -1874
rect 1399 -2062 1445 -2050
rect 1557 -1874 1603 -1862
rect 1557 -2050 1563 -1874
rect 1597 -2050 1603 -1874
rect 1557 -2062 1603 -2050
rect 1715 -1874 1761 -1862
rect 1715 -2050 1721 -1874
rect 1755 -2050 1761 -1874
rect 1715 -2062 1761 -2050
rect 1873 -1874 1919 -1862
rect 1873 -2050 1879 -1874
rect 1913 -2050 1919 -1874
rect 1873 -2062 1919 -2050
rect 2031 -1874 2077 -1862
rect 2031 -2050 2037 -1874
rect 2071 -2050 2077 -1874
rect 2031 -2062 2077 -2050
rect 2189 -1874 2235 -1862
rect 2189 -2050 2195 -1874
rect 2229 -2050 2235 -1874
rect 2189 -2062 2235 -2050
rect -2179 -2109 -2087 -2103
rect -2179 -2143 -2167 -2109
rect -2099 -2143 -2087 -2109
rect -2179 -2149 -2087 -2143
rect -2021 -2109 -1929 -2103
rect -2021 -2143 -2009 -2109
rect -1941 -2143 -1929 -2109
rect -2021 -2149 -1929 -2143
rect -1863 -2109 -1771 -2103
rect -1863 -2143 -1851 -2109
rect -1783 -2143 -1771 -2109
rect -1863 -2149 -1771 -2143
rect -1705 -2109 -1613 -2103
rect -1705 -2143 -1693 -2109
rect -1625 -2143 -1613 -2109
rect -1705 -2149 -1613 -2143
rect -1547 -2109 -1455 -2103
rect -1547 -2143 -1535 -2109
rect -1467 -2143 -1455 -2109
rect -1547 -2149 -1455 -2143
rect -1389 -2109 -1297 -2103
rect -1389 -2143 -1377 -2109
rect -1309 -2143 -1297 -2109
rect -1389 -2149 -1297 -2143
rect -1231 -2109 -1139 -2103
rect -1231 -2143 -1219 -2109
rect -1151 -2143 -1139 -2109
rect -1231 -2149 -1139 -2143
rect -1073 -2109 -981 -2103
rect -1073 -2143 -1061 -2109
rect -993 -2143 -981 -2109
rect -1073 -2149 -981 -2143
rect -915 -2109 -823 -2103
rect -915 -2143 -903 -2109
rect -835 -2143 -823 -2109
rect -915 -2149 -823 -2143
rect -757 -2109 -665 -2103
rect -757 -2143 -745 -2109
rect -677 -2143 -665 -2109
rect -757 -2149 -665 -2143
rect -599 -2109 -507 -2103
rect -599 -2143 -587 -2109
rect -519 -2143 -507 -2109
rect -599 -2149 -507 -2143
rect -441 -2109 -349 -2103
rect -441 -2143 -429 -2109
rect -361 -2143 -349 -2109
rect -441 -2149 -349 -2143
rect -283 -2109 -191 -2103
rect -283 -2143 -271 -2109
rect -203 -2143 -191 -2109
rect -283 -2149 -191 -2143
rect -125 -2109 -33 -2103
rect -125 -2143 -113 -2109
rect -45 -2143 -33 -2109
rect -125 -2149 -33 -2143
rect 33 -2109 125 -2103
rect 33 -2143 45 -2109
rect 113 -2143 125 -2109
rect 33 -2149 125 -2143
rect 191 -2109 283 -2103
rect 191 -2143 203 -2109
rect 271 -2143 283 -2109
rect 191 -2149 283 -2143
rect 349 -2109 441 -2103
rect 349 -2143 361 -2109
rect 429 -2143 441 -2109
rect 349 -2149 441 -2143
rect 507 -2109 599 -2103
rect 507 -2143 519 -2109
rect 587 -2143 599 -2109
rect 507 -2149 599 -2143
rect 665 -2109 757 -2103
rect 665 -2143 677 -2109
rect 745 -2143 757 -2109
rect 665 -2149 757 -2143
rect 823 -2109 915 -2103
rect 823 -2143 835 -2109
rect 903 -2143 915 -2109
rect 823 -2149 915 -2143
rect 981 -2109 1073 -2103
rect 981 -2143 993 -2109
rect 1061 -2143 1073 -2109
rect 981 -2149 1073 -2143
rect 1139 -2109 1231 -2103
rect 1139 -2143 1151 -2109
rect 1219 -2143 1231 -2109
rect 1139 -2149 1231 -2143
rect 1297 -2109 1389 -2103
rect 1297 -2143 1309 -2109
rect 1377 -2143 1389 -2109
rect 1297 -2149 1389 -2143
rect 1455 -2109 1547 -2103
rect 1455 -2143 1467 -2109
rect 1535 -2143 1547 -2109
rect 1455 -2149 1547 -2143
rect 1613 -2109 1705 -2103
rect 1613 -2143 1625 -2109
rect 1693 -2143 1705 -2109
rect 1613 -2149 1705 -2143
rect 1771 -2109 1863 -2103
rect 1771 -2143 1783 -2109
rect 1851 -2143 1863 -2109
rect 1771 -2149 1863 -2143
rect 1929 -2109 2021 -2103
rect 1929 -2143 1941 -2109
rect 2009 -2143 2021 -2109
rect 1929 -2149 2021 -2143
rect 2087 -2109 2179 -2103
rect 2087 -2143 2099 -2109
rect 2167 -2143 2179 -2109
rect 2087 -2149 2179 -2143
<< properties >>
string FIXED_BBOX -2346 -2264 2346 2264
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 10 nf 28 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
