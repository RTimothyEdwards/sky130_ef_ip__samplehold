magic
tech sky130A
magscale 1 2
timestamp 1651948471
<< pwell >>
rect -1632 -1598 1632 1598
<< psubdiff >>
rect -1596 1528 -1500 1562
rect 1500 1528 1596 1562
rect -1596 1466 -1562 1528
rect 1562 1466 1596 1528
rect -1596 -1528 -1562 -1466
rect 1562 -1528 1596 -1466
rect -1596 -1562 -1500 -1528
rect 1500 -1562 1596 -1528
<< psubdiffcont >>
rect -1500 1528 1500 1562
rect -1596 -1466 -1562 1466
rect 1562 -1466 1596 1466
rect -1500 -1562 1500 -1528
<< xpolycontact >>
rect -1466 1000 -1396 1432
rect -1466 -1432 -1396 -1000
rect -1148 1000 -1078 1432
rect -1148 -1432 -1078 -1000
rect -830 1000 -760 1432
rect -830 -1432 -760 -1000
rect -512 1000 -442 1432
rect -512 -1432 -442 -1000
rect -194 1000 -124 1432
rect -194 -1432 -124 -1000
rect 124 1000 194 1432
rect 124 -1432 194 -1000
rect 442 1000 512 1432
rect 442 -1432 512 -1000
rect 760 1000 830 1432
rect 760 -1432 830 -1000
rect 1078 1000 1148 1432
rect 1078 -1432 1148 -1000
rect 1396 1000 1466 1432
rect 1396 -1432 1466 -1000
<< xpolyres >>
rect -1466 -1000 -1396 1000
rect -1148 -1000 -1078 1000
rect -830 -1000 -760 1000
rect -512 -1000 -442 1000
rect -194 -1000 -124 1000
rect 124 -1000 194 1000
rect 442 -1000 512 1000
rect 760 -1000 830 1000
rect 1078 -1000 1148 1000
rect 1396 -1000 1466 1000
<< locali >>
rect -1596 1528 -1500 1562
rect 1500 1528 1596 1562
rect -1596 1466 -1562 1528
rect 1562 1466 1596 1528
rect -1596 -1528 -1562 -1466
rect 1562 -1528 1596 -1466
rect -1596 -1562 -1500 -1528
rect 1500 -1562 1596 -1528
<< viali >>
rect -1450 1017 -1412 1414
rect -1132 1017 -1094 1414
rect -814 1017 -776 1414
rect -496 1017 -458 1414
rect -178 1017 -140 1414
rect 140 1017 178 1414
rect 458 1017 496 1414
rect 776 1017 814 1414
rect 1094 1017 1132 1414
rect 1412 1017 1450 1414
rect -1450 -1414 -1412 -1017
rect -1132 -1414 -1094 -1017
rect -814 -1414 -776 -1017
rect -496 -1414 -458 -1017
rect -178 -1414 -140 -1017
rect 140 -1414 178 -1017
rect 458 -1414 496 -1017
rect 776 -1414 814 -1017
rect 1094 -1414 1132 -1017
rect 1412 -1414 1450 -1017
<< metal1 >>
rect -1456 1414 -1406 1426
rect -1456 1017 -1450 1414
rect -1412 1017 -1406 1414
rect -1456 1005 -1406 1017
rect -1138 1414 -1088 1426
rect -1138 1017 -1132 1414
rect -1094 1017 -1088 1414
rect -1138 1005 -1088 1017
rect -820 1414 -770 1426
rect -820 1017 -814 1414
rect -776 1017 -770 1414
rect -820 1005 -770 1017
rect -502 1414 -452 1426
rect -502 1017 -496 1414
rect -458 1017 -452 1414
rect -502 1005 -452 1017
rect -184 1414 -134 1426
rect -184 1017 -178 1414
rect -140 1017 -134 1414
rect -184 1005 -134 1017
rect 134 1414 184 1426
rect 134 1017 140 1414
rect 178 1017 184 1414
rect 134 1005 184 1017
rect 452 1414 502 1426
rect 452 1017 458 1414
rect 496 1017 502 1414
rect 452 1005 502 1017
rect 770 1414 820 1426
rect 770 1017 776 1414
rect 814 1017 820 1414
rect 770 1005 820 1017
rect 1088 1414 1138 1426
rect 1088 1017 1094 1414
rect 1132 1017 1138 1414
rect 1088 1005 1138 1017
rect 1406 1414 1456 1426
rect 1406 1017 1412 1414
rect 1450 1017 1456 1414
rect 1406 1005 1456 1017
rect -1456 -1017 -1406 -1005
rect -1456 -1414 -1450 -1017
rect -1412 -1414 -1406 -1017
rect -1456 -1426 -1406 -1414
rect -1138 -1017 -1088 -1005
rect -1138 -1414 -1132 -1017
rect -1094 -1414 -1088 -1017
rect -1138 -1426 -1088 -1414
rect -820 -1017 -770 -1005
rect -820 -1414 -814 -1017
rect -776 -1414 -770 -1017
rect -820 -1426 -770 -1414
rect -502 -1017 -452 -1005
rect -502 -1414 -496 -1017
rect -458 -1414 -452 -1017
rect -502 -1426 -452 -1414
rect -184 -1017 -134 -1005
rect -184 -1414 -178 -1017
rect -140 -1414 -134 -1017
rect -184 -1426 -134 -1414
rect 134 -1017 184 -1005
rect 134 -1414 140 -1017
rect 178 -1414 184 -1017
rect 134 -1426 184 -1414
rect 452 -1017 502 -1005
rect 452 -1414 458 -1017
rect 496 -1414 502 -1017
rect 452 -1426 502 -1414
rect 770 -1017 820 -1005
rect 770 -1414 776 -1017
rect 814 -1414 820 -1017
rect 770 -1426 820 -1414
rect 1088 -1017 1138 -1005
rect 1088 -1414 1094 -1017
rect 1132 -1414 1138 -1017
rect 1088 -1426 1138 -1414
rect 1406 -1017 1456 -1005
rect 1406 -1414 1412 -1017
rect 1450 -1414 1456 -1017
rect 1406 -1426 1456 -1414
<< res0p35 >>
rect -1468 -1002 -1394 1002
rect -1150 -1002 -1076 1002
rect -832 -1002 -758 1002
rect -514 -1002 -440 1002
rect -196 -1002 -122 1002
rect 122 -1002 196 1002
rect 440 -1002 514 1002
rect 758 -1002 832 1002
rect 1076 -1002 1150 1002
rect 1394 -1002 1468 1002
<< properties >>
string FIXED_BBOX -1579 -1545 1579 1545
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 10 m 1 nx 10 wmin 0.350 lmin 0.50 rho 2000 val 58.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
