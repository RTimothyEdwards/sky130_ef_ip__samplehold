magic
tech sky130A
magscale 1 2
timestamp 1718228984
<< error_s >>
rect 10732 10710 10835 10726
rect 11721 10710 12149 10726
rect 10704 10682 10835 10698
rect 11721 10682 12177 10698
rect 2512 10548 3512 10621
rect 4440 10548 5440 10621
rect 2512 9621 2599 10548
rect 5353 9621 5440 10548
rect 5898 10548 6898 10621
rect 7826 10548 8826 10621
rect 5898 9621 5985 10548
rect 8739 9621 8826 10548
rect 9284 10548 10284 10621
rect 11212 10548 12212 10621
rect 9284 9621 9371 10548
rect 10983 10325 11005 10401
rect 11011 10353 11033 10429
rect 10983 10191 11008 10325
rect 11011 10163 11036 10353
rect 11402 10251 11403 10441
rect 11430 10279 11431 10413
rect 10983 9889 11005 9965
rect 10983 9755 11008 9889
rect 10983 9453 11005 9529
rect 2512 8332 2599 9332
rect 5353 8332 5440 9332
rect 5898 8332 5985 9332
rect 8739 8332 8826 9332
rect 9284 8332 9371 9332
rect 10983 9319 11008 9453
rect 11011 9266 11403 10153
rect 11430 9930 11431 9977
rect 11424 9849 11431 9930
rect 11430 9843 11431 9849
rect 12125 9621 12212 10548
rect 12670 10548 13670 10621
rect 14598 10548 15598 10621
rect 12670 9621 12757 10548
rect 15511 9621 15598 10548
rect 16056 10548 17056 10621
rect 17984 10548 18984 10621
rect 16056 9621 16143 10548
rect 18897 9621 18984 10548
rect 11430 9494 11431 9541
rect 11424 9413 11431 9494
rect 11430 9407 11431 9413
rect 10983 9017 11005 9093
rect 11011 9045 11033 9121
rect 11402 9058 11403 9133
rect 11430 9058 11431 9105
rect 10983 8883 11008 9017
rect 11011 8855 11036 9045
rect 11396 8949 11403 9058
rect 11424 8977 11431 9058
rect 11430 8971 11431 8977
rect 11402 8943 11403 8949
rect 10983 8581 11005 8657
rect 11011 8609 11033 8685
rect 11402 8622 11403 8697
rect 11430 8622 11431 8669
rect 10983 8447 11008 8581
rect 11011 8419 11036 8609
rect 11396 8513 11403 8622
rect 11424 8541 11431 8622
rect 11430 8535 11431 8541
rect 11402 8507 11403 8513
rect 12125 8332 12212 9332
rect 12670 8332 12757 9332
rect 15511 8332 15598 9332
rect 16056 8332 16143 9332
rect 18897 8332 18984 9332
rect 10983 8145 11005 8221
rect 11011 8173 11033 8249
rect 11402 8186 11403 8261
rect 11430 8186 11431 8233
rect 2512 7043 2599 8043
rect 5353 7043 5440 8043
rect 5898 7043 5985 8043
rect 8739 7043 8826 8043
rect 9284 7043 9371 8043
rect 10983 8011 11008 8145
rect 11011 7983 11036 8173
rect 11396 8077 11403 8186
rect 11424 8105 11431 8186
rect 11430 8099 11431 8105
rect 11402 8071 11403 8077
rect 10983 7709 11005 7785
rect 11011 7737 11033 7813
rect 11402 7750 11403 7825
rect 11430 7750 11431 7797
rect 10983 7575 11008 7709
rect 11011 7547 11036 7737
rect 11396 7641 11403 7750
rect 11424 7669 11431 7750
rect 11430 7663 11431 7669
rect 11402 7635 11403 7641
rect 10983 7273 11005 7349
rect 11011 7301 11033 7377
rect 11402 7314 11403 7389
rect 11430 7314 11431 7361
rect 10983 7139 11008 7273
rect 11011 7111 11036 7301
rect 11396 7205 11403 7314
rect 11424 7233 11431 7314
rect 11430 7227 11431 7233
rect 11402 7199 11403 7205
rect 12125 7043 12212 8043
rect 12670 7043 12757 8043
rect 15511 7043 15598 8043
rect 16056 7043 16143 8043
rect 18897 7043 18984 8043
rect 10983 6837 11005 6913
rect 11011 6865 11033 6941
rect 11402 6878 11403 6953
rect 11430 6878 11431 6925
rect 2512 5754 2599 6754
rect 5353 5754 5440 6754
rect 5898 5754 5985 6754
rect 8739 5754 8826 6754
rect 9284 5754 9371 6754
rect 10983 6703 11008 6837
rect 11011 6675 11036 6865
rect 11396 6769 11403 6878
rect 11424 6797 11431 6878
rect 11430 6791 11431 6797
rect 11402 6763 11403 6769
rect 10983 6401 11005 6477
rect 11011 6429 11033 6505
rect 11402 6442 11403 6517
rect 11430 6442 11431 6489
rect 10983 6267 11008 6401
rect 11011 6327 11036 6429
rect 11272 6327 11324 6395
rect 11396 6333 11403 6442
rect 11424 6361 11431 6442
rect 11430 6355 11431 6361
rect 11402 6327 11403 6333
rect 11011 6239 11387 6327
rect 11029 6069 11387 6239
rect 10983 5965 11005 6041
rect 11011 5969 11387 6069
rect 11402 6006 11403 6081
rect 11430 6006 11431 6053
rect 10983 5921 11008 5965
rect 11011 5949 11036 5969
rect 11114 5925 11166 5969
rect 11396 5897 11403 6006
rect 11424 5925 11431 6006
rect 12125 5754 12212 6754
rect 12353 5813 12368 5842
rect 12381 5841 12396 5870
rect 12670 5754 12757 6754
rect 15511 5754 15598 6754
rect 16056 5754 16143 6754
rect 18897 5754 18984 6754
rect 2512 4465 2599 5465
rect 5353 4465 5440 5465
rect 5898 4465 5985 5465
rect 8739 4465 8826 5465
rect 9284 4465 9371 5465
rect 11396 5461 11403 5570
rect 11424 5489 11431 5570
rect 12350 5488 12368 5645
rect 12378 5483 12396 5617
rect 11028 5197 11386 5340
rect 12125 5224 12212 5465
rect 12381 5460 12396 5483
rect 11550 5215 11676 5224
rect 11550 5210 11581 5215
rect 11647 5210 11676 5215
rect 11708 5215 11834 5224
rect 11708 5210 11739 5215
rect 11805 5210 11834 5215
rect 11866 5215 11992 5224
rect 11866 5210 11897 5215
rect 11963 5210 11992 5215
rect 12024 5215 12212 5224
rect 12024 5210 12055 5215
rect 12121 5210 12212 5215
rect 10983 5093 11005 5169
rect 10983 4959 11008 5093
rect 11011 4982 11386 5197
rect 11402 5134 11403 5209
rect 12125 5196 12212 5210
rect 11550 5187 11676 5196
rect 11550 5182 11609 5187
rect 11619 5182 11676 5187
rect 11708 5187 11834 5196
rect 11708 5182 11767 5187
rect 11777 5182 11834 5187
rect 11866 5187 11992 5196
rect 11866 5182 11925 5187
rect 11935 5182 11992 5187
rect 12024 5187 12212 5196
rect 12024 5182 12083 5187
rect 12093 5182 12212 5187
rect 11430 5134 11431 5181
rect 11396 5025 11403 5134
rect 11424 5053 11431 5134
rect 11430 5047 11431 5053
rect 11402 5019 11403 5025
rect 11011 4931 11036 4982
rect 11272 4965 11324 4982
rect 11721 4941 11746 4996
rect 11749 4969 11774 4996
rect 11847 4820 11866 4879
rect 11875 4820 11894 4851
rect 10983 4657 11005 4733
rect 11011 4685 11033 4761
rect 11402 4698 11403 4773
rect 11430 4698 11431 4745
rect 10983 4523 11008 4657
rect 11011 4495 11036 4685
rect 11396 4589 11403 4698
rect 11424 4617 11431 4698
rect 11430 4611 11431 4617
rect 11402 4583 11403 4589
rect 11721 4505 11746 4611
rect 11749 4533 11774 4611
rect 11847 4492 11866 4774
rect 11875 4492 11894 4774
rect 11964 4492 11987 4651
rect 11992 4492 12015 4651
rect 12125 4465 12212 5182
rect 12670 4465 12757 5465
rect 15511 4465 15598 5465
rect 16056 4465 16143 5465
rect 18897 4465 18984 5465
rect 11011 4368 11403 4451
rect 9885 4306 13033 4368
rect 2512 3176 2599 4176
rect 5353 3176 5440 4176
rect 5898 3176 5985 4176
rect 8739 3176 8826 4176
rect 9284 3176 9371 4176
rect 10983 4074 11005 4129
rect 11011 4074 11403 4306
rect 10976 4050 11403 4074
rect 10983 4046 11008 4050
rect 11011 4046 11036 4050
rect 10950 4022 11036 4046
rect 10983 3918 11008 4022
rect 11011 3890 11036 4022
rect 11114 4012 11166 4050
rect 11266 4022 11330 4046
rect 11402 3978 11403 4050
rect 11430 4006 11431 4140
rect 11554 4050 11674 4074
rect 11582 4022 11646 4046
rect 11721 3901 11746 4006
rect 11749 3929 11774 4006
rect 11847 3888 11866 4170
rect 11875 4074 11894 4170
rect 11964 4074 11987 4170
rect 11870 4050 11990 4074
rect 11875 3888 11894 4050
rect 11898 4022 11962 4046
rect 11964 3888 11987 4050
rect 11992 3888 12015 4170
rect 10710 3114 10732 3292
rect 10738 3142 10760 3264
rect 11518 3227 11537 3361
rect 11518 3148 11536 3227
rect 11546 3199 11565 3389
rect 11847 3227 11853 3361
rect 10711 3028 10732 3114
rect 10739 3028 10760 3142
rect 11546 3120 11564 3199
rect 11847 3148 11852 3227
rect 11875 3199 11881 3389
rect 11875 3120 11880 3199
rect 12125 3176 12212 4176
rect 12670 3176 12757 4176
rect 15511 3176 15598 4176
rect 16056 3176 16143 4176
rect 18897 3176 18984 4176
rect 2512 1887 2599 2887
rect 3648 1925 3657 2298
rect 3676 1897 3685 2326
rect 5353 1887 5440 2887
rect 5898 1887 5985 2887
rect 8739 1887 8826 2887
rect 9284 1887 9371 2887
rect 11981 2575 11987 2793
rect 12009 2575 12015 2793
rect 11867 2378 11933 2382
rect 11868 2376 11932 2378
rect 10896 2372 10921 2374
rect 11022 2299 11074 2301
rect 11011 1920 11403 2289
rect 11981 2265 11987 2529
rect 12009 2265 12015 2529
rect 9971 1868 11985 1920
rect 12125 1887 12212 2887
rect 12670 1887 12757 2887
rect 15511 1887 15598 2887
rect 16056 1887 16143 2887
rect 18897 1887 18984 2887
rect 2512 598 2599 1598
rect 5353 598 5440 1598
rect 5898 598 5985 1598
rect 8739 598 8826 1598
rect 9284 598 9371 1598
rect 10896 1577 10923 1657
rect 10983 1469 10984 1692
rect 10896 1107 10952 1119
rect 11011 1096 11403 1868
rect 11744 1273 11746 1730
rect 11772 1301 11774 1702
rect 11921 1577 11942 1595
rect 11936 1521 11998 1539
rect 11957 1393 11977 1426
rect 12125 1096 12212 1598
rect 9799 1033 12566 1096
rect 11011 660 11403 1033
rect 12125 598 12212 1033
rect 12670 598 12757 1598
rect 15511 598 15598 1598
rect 16056 598 16143 1598
rect 18897 598 18984 1598
rect 11885 440 12206 483
rect 9652 379 13186 440
rect 11885 370 12206 379
<< locali >>
rect 392 8914 616 9238
rect 940 9208 2054 9238
rect 940 8946 1166 9208
rect 2008 8946 2054 9208
rect 940 8914 2054 8946
rect 392 8734 426 8914
rect 2020 8732 2054 8914
rect 722 8622 830 8646
rect 722 8262 744 8622
rect 814 8262 830 8622
rect 722 8214 830 8262
rect 1692 6610 1778 6648
rect 1428 6600 1778 6610
rect 1428 6536 1440 6600
rect 1764 6536 1778 6600
rect 1428 6524 1778 6536
<< viali >>
rect 1166 8946 2008 9208
rect 744 8262 814 8622
rect 1440 6536 1764 6600
<< metal1 >>
rect 11011 11170 11403 11182
rect 11011 10890 11023 11170
rect 11389 10890 11403 11170
rect 11011 10153 11403 10890
rect 0 9612 1070 9952
rect 0 9040 200 9101
rect 0 8950 815 9040
rect 0 8901 200 8950
rect 743 8632 815 8950
rect 1013 8655 1070 9612
rect 1118 9208 2060 9238
rect 1118 8946 1166 9208
rect 2008 8946 2060 9208
rect 1118 8914 2060 8946
rect 1912 8702 1986 8914
rect 2014 8738 2060 8914
rect 2014 8702 2020 8738
rect 2054 8702 2060 8738
rect 732 8622 826 8632
rect 732 8262 744 8622
rect 814 8262 826 8622
rect 732 8246 826 8262
rect 386 6474 432 6652
rect 460 6474 534 6652
rect 0 6462 1040 6474
rect 0 6166 814 6462
rect 1026 6166 1040 6462
rect 0 6152 1040 6166
rect 1098 6082 1172 6700
rect 1200 6082 1246 6646
rect 1274 6082 1348 6700
rect 1428 6600 1778 6610
rect 1428 6536 1440 6600
rect 1764 6536 1778 6600
rect 1428 6524 1778 6536
rect 1912 6476 1986 6640
rect 2014 6476 2060 6640
rect 1406 6464 2060 6476
rect 1406 6168 1422 6464
rect 1616 6168 2060 6464
rect 1406 6152 2060 6168
rect 11011 6327 11403 9266
rect 1098 6015 1348 6082
rect 0 5284 2515 6015
rect 3391 5284 3424 6015
rect 11011 5969 11029 6327
rect 11387 5969 11403 6327
rect 11011 5949 11403 5969
rect 10725 5488 12368 5842
rect 11011 5340 11403 5360
rect 0 4986 3717 5186
rect 11011 4982 11028 5340
rect 11386 4982 11403 5340
rect 0 4641 1888 4841
rect 2381 4641 3717 4841
rect 11011 4451 11403 4982
rect 2404 2443 2515 2719
rect 3391 2443 3517 2719
rect 2924 1925 3657 2298
rect 11011 2289 11403 4050
rect 2416 1647 2693 1847
rect 2493 1595 2693 1647
rect 2493 1427 2693 1436
rect 2924 1287 3506 1925
rect 2924 941 2942 1287
rect 2402 726 2942 941
rect 3484 726 3506 1287
rect 2402 706 3506 726
rect 11011 627 11403 660
rect 11546 4996 12150 5196
rect 11546 281 11746 4996
rect 11875 4651 12150 4851
rect 11875 483 11987 4651
rect 19130 4570 19469 4770
rect 11875 370 11885 483
rect 12206 370 12216 483
rect 2478 248 3021 281
rect 2478 -80 2519 248
rect 2985 -80 3021 248
rect 2478 -114 3021 -80
rect 11278 248 11821 281
rect 11278 -80 11319 248
rect 11785 -80 11821 248
rect 11278 -114 11821 -80
<< via1 >>
rect 11023 10890 11389 11170
rect 11011 9266 11403 10153
rect 814 6166 1026 6462
rect 1440 6536 1764 6600
rect 1422 6168 1616 6464
rect 2515 5284 3391 6015
rect 11029 5969 11387 6327
rect 11028 4982 11386 5340
rect 1888 4641 2381 4841
rect 11011 4050 11403 4451
rect 2515 2443 3391 2719
rect 2493 1436 2693 1595
rect 872 718 1589 929
rect 2942 726 3484 1287
rect 11011 660 11403 2289
rect 11885 370 12206 483
rect 2519 -80 2985 248
rect 11319 -80 11785 248
<< metal2 >>
rect 11011 11170 11403 11182
rect 2515 10932 3391 11027
rect 2515 10710 3685 10932
rect 10732 10756 10958 10932
rect 11011 10890 11023 11170
rect 11389 10890 11403 11170
rect 11011 10836 11403 10890
rect 11477 10756 12149 10942
rect 10732 10710 12149 10756
rect 1428 6600 1778 6610
rect 1428 6536 1440 6600
rect 1764 6536 1778 6600
rect 1428 6524 1778 6536
rect 798 6464 1630 6474
rect 798 6462 1422 6464
rect 798 6166 814 6462
rect 1026 6168 1422 6462
rect 1616 6168 1630 6464
rect 1026 6166 1630 6168
rect 798 6152 1630 6166
rect 1692 3414 1778 6524
rect 2515 6015 3391 10710
rect 10835 10479 11721 10710
rect 11011 10153 11403 10231
rect 11011 6327 11403 9266
rect 11011 5969 11029 6327
rect 11387 5969 11403 6327
rect 3391 5573 3685 5842
rect 1871 4641 1888 4841
rect 2381 4641 2394 4841
rect 856 929 1605 940
rect 856 718 872 929
rect 1589 718 1605 929
rect 856 706 1605 718
rect 2300 464 2394 4641
rect 2515 2719 3391 5284
rect 11011 5340 11403 5969
rect 11011 4982 11028 5340
rect 11386 4982 11403 5340
rect 2515 2403 3391 2443
rect 10573 1595 10732 4882
rect 11011 4451 11403 4982
rect 10976 4050 11011 4451
rect 11403 4050 12119 4451
rect 2484 1436 2493 1595
rect 2693 1436 10732 1595
rect 10952 2289 12119 2326
rect 2924 1287 3506 1305
rect 2924 726 2942 1287
rect 3484 803 3506 1287
rect 10952 803 11011 2289
rect 3484 726 11011 803
rect 2924 660 11011 726
rect 11403 1934 12119 2289
rect 11403 803 11921 1934
rect 11403 660 19235 803
rect 2924 578 19235 660
rect 11875 464 11885 483
rect 2300 370 11885 464
rect 12206 370 12216 483
rect 2478 248 3021 281
rect 2478 -80 2519 248
rect 2985 -80 3021 248
rect 2478 -114 3021 -80
rect 11278 248 11821 281
rect 11278 -80 11319 248
rect 11785 -80 11821 248
rect 11278 -114 11821 -80
<< via2 >>
rect 11023 10890 11389 11170
rect 357 1087 508 2307
rect 872 718 1589 929
rect 2519 -80 2985 248
rect 11319 -80 11785 248
<< metal3 >>
rect 11011 11170 11403 11182
rect 11011 10890 11023 11170
rect 11389 10890 11403 11170
rect 11011 10879 11403 10890
rect 337 2307 522 2321
rect 337 1087 357 2307
rect 508 1087 522 2307
rect 337 191 522 1087
rect 856 929 1605 940
rect 856 718 872 929
rect 1589 718 1605 929
rect 856 706 1605 718
rect 2478 248 3021 281
rect 2478 191 2519 248
rect 337 6 2519 191
rect 2478 -80 2519 6
rect 2985 -80 3021 248
rect 2478 -114 3021 -80
rect 11278 248 11821 281
rect 11278 -80 11319 248
rect 11785 -80 11821 248
rect 11278 -114 11821 -80
<< via3 >>
rect 11023 10890 11389 11170
rect 872 718 1589 929
rect 2519 -80 2985 248
rect 11319 -80 11785 248
<< metal4 >>
rect 0 11182 1039 11183
rect 0 10817 2236 11182
rect 0 10191 1606 10817
rect 857 929 1606 10191
rect 857 718 872 929
rect 1589 718 1606 929
rect 857 637 1606 718
rect 2478 248 3021 281
rect 2478 -80 2519 248
rect 2985 -80 3021 248
rect 2478 -114 3021 -80
rect 11278 248 11821 281
rect 11278 -80 11319 248
rect 11785 -80 11821 248
rect 11278 -114 11821 -80
<< via4 >>
rect 2519 -80 2985 248
rect 11319 -80 11785 248
<< metal5 >>
rect 2478 248 3021 281
rect 2478 -80 2519 248
rect 2985 -80 3021 248
rect 2478 -114 3021 -80
rect 11278 248 11871 281
rect 11278 -80 11319 248
rect 11785 -80 11871 248
rect 11278 -114 11871 -80
use hold_cap_array  hold_cap_array_0
timestamp 1652200182
transform 1 0 218 0 1 26439
box 1997 -26553 19047 -15257
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_0 paramcells
timestamp 1652928066
transform 1 0 778 0 1 9076
box -198 -198 198 198
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 0 1 409 -1 0 8738
box -66 -43 2178 1671
use balanced_switch  x1
timestamp 1718228984
transform -1 0 2730 0 1 2811
box 301 -2311 2543 1830
use follower_amp  x2
timestamp 1718228984
transform 1 0 3676 0 1 -174
box 0 0 4377 11129
use follower_amp  x3
timestamp 1718228984
transform 1 0 9246 0 1 -84
box 0 0 4377 11129
<< labels >>
flabel metal1 0 5284 200 6015 0 FreeSans 320 0 0 0 vdd
port 2 nsew
flabel metal1 0 8901 200 9101 0 FreeSans 256 0 0 0 hold
port 3 nsew
flabel metal1 0 9612 804 9952 0 FreeSans 1600 0 0 0 dvdd
port 6 nsew
flabel metal1 0 6152 788 6474 0 FreeSans 1600 0 0 0 dvss
port 7 nsew
flabel metal4 0 10191 1039 11183 0 FreeSans 1600 0 0 0 vss
port 5 nsew
flabel metal1 19269 4570 19469 4770 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 0 4986 200 5186 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal1 0 4641 200 4841 0 FreeSans 320 0 0 0 ena
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 19469 11297
<< end >>
