magic
tech sky130A
magscale 1 2
timestamp 1651944383
<< error_p >>
rect -96 333 -62 353
rect -50 333 50 391
rect 62 333 96 353
rect -108 331 108 333
rect -133 307 -108 331
rect -96 327 -62 331
rect -50 327 -25 331
rect 25 327 50 331
rect 62 327 96 331
rect -104 307 104 327
rect 108 307 133 331
rect -133 306 133 307
rect -130 298 130 306
rect -133 285 133 298
rect -133 273 -108 285
rect -104 273 104 285
rect 108 273 133 285
rect -296 100 -263 273
rect -242 138 -209 273
rect -96 197 -62 228
rect -50 213 50 273
rect -50 197 -49 198
rect -45 197 0 213
rect 49 197 50 198
rect 62 197 96 228
rect 108 197 154 255
rect -180 181 2 197
rect 50 191 180 197
rect -134 147 -129 181
rect -113 171 -49 181
rect -108 157 -49 171
rect -113 147 -49 157
rect -45 147 2 181
rect 35 181 180 191
rect 35 147 45 181
rect 50 147 113 181
rect 129 147 134 181
rect -242 100 -196 138
rect -180 137 -35 147
rect 35 137 180 147
rect 209 138 242 273
rect -180 101 -108 137
rect -96 101 -36 137
rect 62 101 180 137
rect -180 100 -107 101
rect -97 100 -36 101
rect 61 100 180 101
rect 196 100 242 138
rect 263 100 296 273
rect -327 -100 -321 100
rect -296 -100 -196 100
rect -187 75 -159 100
rect -187 -75 -184 75
rect -175 -75 -162 75
rect -134 74 -127 100
rect -109 99 -108 100
rect -96 99 -95 100
rect -63 99 -62 100
rect 62 99 63 100
rect 95 99 96 100
rect 108 99 109 100
rect -28 88 28 99
rect -129 -74 -127 74
rect -187 -100 -159 -75
rect -134 -100 -127 -74
rect -17 -77 -6 88
rect 17 -77 28 88
rect -17 -88 28 -77
rect 127 74 134 100
rect 159 75 184 100
rect 127 -74 129 74
rect -109 -100 -108 -99
rect -96 -100 -95 -99
rect -63 -100 -62 -99
rect 62 -100 63 -99
rect 95 -100 96 -99
rect 108 -100 109 -99
rect 127 -100 134 -74
rect 162 -75 175 75
rect 159 -100 184 -75
rect 196 -100 296 100
rect 321 -100 327 100
rect -296 -273 -263 -100
rect -242 -138 -196 -100
rect -180 -101 -107 -100
rect -97 -101 2 -100
rect 61 -101 180 -100
rect -180 -137 -108 -101
rect -96 -137 2 -101
rect 62 -137 180 -101
rect -242 -273 -209 -138
rect -180 -147 2 -137
rect -134 -181 -129 -147
rect -113 -157 -49 -147
rect -108 -171 -49 -157
rect -113 -181 -49 -171
rect -45 -181 2 -147
rect 35 -147 180 -137
rect 196 -138 242 -100
rect 35 -181 45 -147
rect 50 -181 113 -147
rect 129 -181 134 -147
rect -180 -191 -35 -181
rect 35 -191 180 -181
rect -180 -197 -36 -191
rect 50 -197 180 -191
rect -50 -198 -49 -197
rect 49 -198 50 -197
rect -96 -271 -62 -251
rect -50 -271 50 -213
rect 62 -271 96 -251
rect -108 -273 108 -271
rect 209 -273 242 -138
rect 263 -273 296 -100
rect -133 -297 -108 -273
rect -96 -277 -62 -273
rect -50 -277 -25 -273
rect 25 -277 50 -273
rect 62 -277 96 -273
rect -104 -297 104 -277
rect 108 -297 133 -273
rect -133 -298 133 -297
rect -130 -306 130 -298
rect -133 -319 133 -306
rect -133 -331 -108 -319
rect -104 -331 104 -319
rect 108 -331 133 -319
rect -50 -391 50 -331
<< nwell >>
rect -308 397 308 797
rect -387 -397 387 397
rect -308 -797 308 -397
<< mvpmos >>
rect -50 331 50 500
rect -50 197 50 273
rect -108 181 -96 197
rect -62 181 62 197
rect 96 181 108 197
rect -45 147 45 181
rect -108 100 -96 147
rect -62 100 62 147
rect 96 100 108 147
rect -129 88 129 100
rect -129 -88 -17 88
rect 17 -88 129 88
rect -129 -100 129 -88
rect -108 -147 -96 -100
rect -62 -147 62 -100
rect 96 -147 108 -100
rect -45 -181 45 -147
rect -108 -197 -96 -181
rect -62 -197 62 -181
rect 96 -197 108 -181
rect -50 -273 50 -197
rect -50 -500 50 -331
<< mvpdiff >>
rect -108 488 -50 500
rect -108 331 -96 488
rect -62 331 -50 488
rect 50 488 108 500
rect 50 331 62 488
rect 96 331 108 488
rect -108 197 -96 273
rect -62 197 -50 273
rect 50 197 62 273
rect 96 197 108 273
rect -187 88 -129 100
rect 129 88 187 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect 129 -88 141 88
rect 175 -88 187 88
rect -187 -100 -129 -88
rect 129 -100 187 -88
rect -108 -273 -96 -197
rect -62 -273 -50 -197
rect 50 -273 62 -197
rect 96 -273 108 -197
rect -108 -488 -96 -331
rect -62 -488 -50 -331
rect -108 -500 -50 -488
rect 50 -488 62 -331
rect 96 -488 108 -331
rect 50 -500 108 -488
<< mvpdiffc >>
rect -96 331 -62 488
rect 62 331 96 488
rect -96 197 -62 273
rect 62 197 96 273
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect -96 -273 -62 -197
rect 62 -273 96 -197
rect -96 -488 -62 -331
rect 62 -488 96 -331
<< mvnsubdiff >>
rect -242 719 242 731
rect -242 685 -134 719
rect 134 685 242 719
rect -242 673 242 685
rect -242 623 -184 673
rect -242 331 -230 623
rect -321 273 -230 331
rect -196 331 -184 623
rect 184 623 242 673
rect 184 331 196 623
rect -196 319 196 331
rect 230 331 242 623
rect -321 223 -263 273
rect -321 -223 -309 223
rect -275 -223 -263 223
rect -321 -273 -263 -223
rect -242 -273 -230 273
rect -321 -331 -230 -273
rect -196 273 196 285
rect -196 100 -184 273
rect 184 100 196 273
rect -196 -100 -187 100
rect 187 -100 196 100
rect -196 -273 -184 -100
rect 184 -273 196 -100
rect -196 -285 196 -273
rect 230 273 321 331
rect 230 -273 242 273
rect 263 223 321 273
rect 263 -223 275 223
rect 309 -223 321 223
rect 263 -273 321 -223
rect -242 -623 -230 -331
rect -196 -331 196 -319
rect -196 -623 -184 -331
rect -242 -673 -184 -623
rect 184 -623 196 -331
rect 230 -331 321 -273
rect 230 -623 242 -331
rect 184 -673 242 -623
rect -242 -685 242 -673
rect -242 -719 -134 -685
rect 134 -719 242 -685
rect -242 -731 242 -719
<< mvnsubdiffcont >>
rect -134 685 134 719
rect -230 319 -196 623
rect 196 319 230 623
rect -230 285 230 319
rect -309 -223 -275 223
rect -230 -285 -196 285
rect 196 -285 230 285
rect 275 -223 309 223
rect -230 -319 230 -285
rect -230 -623 -196 -319
rect 196 -623 230 -319
rect -134 -719 134 -685
<< poly >>
rect -50 581 50 597
rect -50 547 -34 581
rect 34 547 50 581
rect -50 500 50 547
rect -129 181 -108 197
rect -96 181 -62 197
rect 62 181 96 197
rect 108 181 129 197
rect -129 147 -113 181
rect 113 147 129 181
rect -129 100 -108 147
rect -96 100 -62 147
rect 62 100 96 147
rect 108 100 129 147
rect -129 -147 -108 -100
rect -96 -147 -62 -100
rect 62 -147 96 -100
rect 108 -147 129 -100
rect -129 -181 -113 -147
rect 113 -181 129 -147
rect -129 -197 -108 -181
rect -96 -197 -62 -181
rect 62 -197 96 -181
rect 108 -197 129 -181
rect -50 -547 50 -500
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -50 -597 50 -581
<< polycont >>
rect -34 547 34 581
rect -113 147 -45 181
rect 45 147 113 181
rect -113 -181 -45 -147
rect 45 -181 113 -147
rect -34 -581 34 -547
<< locali >>
rect -230 685 -134 719
rect 134 685 230 719
rect -230 623 -196 685
rect 196 623 230 685
rect -50 547 -34 581
rect 34 547 50 581
rect -96 488 -62 504
rect 62 488 96 504
rect -309 285 -230 319
rect 230 285 309 319
rect -309 223 -275 285
rect -309 -285 -275 -223
rect -129 147 -113 181
rect -45 147 -29 181
rect 29 147 45 181
rect 113 147 129 181
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 275 223 309 285
rect 275 -285 309 -223
rect -309 -319 -230 -285
rect 230 -319 309 -285
rect -96 -504 -62 -488
rect 62 -504 96 -488
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -230 -685 -196 -623
rect 196 -685 230 -623
rect -230 -719 -134 -685
rect 134 -719 230 -685
<< viali >>
rect -34 547 34 581
rect -96 331 -62 488
rect -96 319 -62 331
rect 62 331 96 488
rect 62 319 96 331
rect -96 285 -62 319
rect 62 285 96 319
rect -96 273 -62 285
rect -96 197 -62 273
rect -96 181 -62 197
rect 62 273 96 285
rect 62 197 96 273
rect 62 181 96 197
rect -113 147 -45 181
rect 45 147 113 181
rect -175 -88 -141 88
rect -96 -147 -62 147
rect -17 -88 17 88
rect 62 -147 96 147
rect 141 -88 175 88
rect -113 -181 -45 -147
rect 45 -181 113 -147
rect -96 -197 -62 -181
rect -96 -273 -62 -197
rect -96 -285 -62 -273
rect 62 -197 96 -181
rect 62 -273 96 -197
rect 62 -285 96 -273
rect -96 -319 -62 -285
rect 62 -319 96 -285
rect -96 -331 -62 -319
rect -96 -488 -62 -331
rect 62 -331 96 -319
rect 62 -488 96 -331
rect -34 -581 34 -547
<< metal1 >>
rect -46 581 46 587
rect -46 547 -34 581
rect 34 547 46 581
rect -46 541 46 547
rect -102 488 -56 500
rect -102 187 -96 488
rect -125 181 -96 187
rect -62 187 -56 488
rect 56 488 102 500
rect 56 187 62 488
rect -62 181 -33 187
rect -125 147 -113 181
rect -45 147 -33 181
rect -125 141 -96 147
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -102 -141 -96 141
rect -125 -147 -96 -141
rect -62 141 -33 147
rect 33 181 62 187
rect 96 187 102 488
rect 96 181 125 187
rect 33 147 45 181
rect 113 147 125 181
rect 33 141 62 147
rect -62 -141 -56 141
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 56 -141 62 141
rect -62 -147 -33 -141
rect -125 -181 -113 -147
rect -45 -181 -33 -147
rect -125 -187 -96 -181
rect -102 -488 -96 -187
rect -62 -187 -33 -181
rect 33 -147 62 -141
rect 96 141 125 147
rect 96 -141 102 141
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect 96 -147 125 -141
rect 33 -181 45 -147
rect 113 -181 125 -147
rect 33 -187 62 -181
rect -62 -488 -56 -187
rect -102 -500 -56 -488
rect 56 -488 62 -187
rect 96 -187 125 -181
rect 96 -488 102 -187
rect 56 -500 102 -488
rect -46 -547 46 -541
rect -46 -581 -34 -547
rect 34 -581 46 -547
rect -46 -587 46 -581
<< properties >>
string FIXED_BBOX -292 -302 292 302
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
