magic
tech sky130A
magscale 1 2
timestamp 1719257891
<< dnwell >>
rect 410 -3000 2434 1930
<< nwell >>
rect 301 1724 2543 2130
rect 301 782 616 1724
rect 2228 782 2543 1724
rect 301 673 2543 782
rect 301 -2794 616 673
rect 1957 -297 2543 673
rect 2228 -2794 2543 -297
rect 301 -3111 2543 -2794
<< mvnsubdiff >>
rect 367 2044 2477 2064
rect 367 2010 447 2044
rect 2397 2010 2477 2044
rect 367 1990 2477 2010
rect 367 1984 441 1990
rect 367 -2963 387 1984
rect 421 -2963 441 1984
rect 367 -2969 441 -2963
rect 2403 1984 2477 1990
rect 2403 -2963 2423 1984
rect 2457 -2963 2477 1984
rect 2403 -2969 2477 -2963
rect 367 -2989 2477 -2969
rect 367 -3023 447 -2989
rect 2397 -3023 2477 -2989
rect 367 -3043 2477 -3023
<< mvnsubdiffcont >>
rect 447 2010 2397 2044
rect 387 -2963 421 1984
rect 2423 -2963 2457 1984
rect 447 -3023 2397 -2989
<< locali >>
rect 387 2010 447 2044
rect 2397 2010 2457 2044
rect 387 1984 2457 2010
rect 421 1921 2423 1984
rect 421 782 571 1921
rect 616 856 768 1676
rect 1169 1655 1343 1677
rect 1169 974 1221 1655
rect 1297 974 1343 1655
rect 1169 856 1343 974
rect 1753 1657 2255 1677
rect 1753 976 1802 1657
rect 1878 1147 2255 1657
rect 1878 976 1927 1147
rect 1753 856 1927 976
rect 2164 856 2255 1147
rect 2325 782 2423 1921
rect 421 642 2423 782
rect 421 -158 712 642
rect 1870 -158 2423 642
rect 421 -185 2423 -158
rect 421 -358 537 -185
rect 2337 -358 2423 -185
rect 421 -374 2423 -358
rect 421 -1694 712 -374
rect 2140 -1694 2423 -374
rect 421 -1788 2423 -1694
rect 421 -2628 528 -1788
rect 599 -1955 2235 -1866
rect 599 -2670 714 -1955
rect 2120 -2670 2235 -1955
rect 2302 -2621 2423 -1788
rect 471 -2711 2378 -2670
rect 471 -2881 582 -2711
rect 2327 -2881 2378 -2711
rect 471 -2943 2378 -2881
rect 387 -2989 421 -2963
rect 2423 -2989 2457 -2963
rect 387 -3023 447 -2989
rect 2397 -3023 2457 -2989
<< viali >>
rect 1221 974 1297 1655
rect 1802 976 1878 1657
rect 537 -358 2337 -185
rect 582 -2881 2327 -2711
<< metal1 >>
rect 393 1841 2463 1863
rect 393 1622 544 1841
rect 842 1657 2463 1841
rect 842 1655 1802 1657
rect 842 1622 1221 1655
rect 393 1606 1221 1622
rect 824 1064 888 1606
rect 340 919 540 990
rect 943 919 980 1531
rect 340 867 894 919
rect 972 867 980 919
rect 340 790 540 867
rect 943 701 980 867
rect 1052 802 1101 1472
rect 1211 974 1221 1606
rect 1297 1606 1802 1655
rect 1297 974 1308 1606
rect 1406 1060 1470 1606
rect 1211 959 1308 974
rect 1534 802 1571 1532
rect 1052 753 1571 802
rect 909 664 1099 701
rect 909 500 946 664
rect 1062 500 1099 664
rect 793 438 866 453
rect 793 -46 803 438
rect 857 -46 866 438
rect 793 -59 866 -46
rect 964 -92 1036 456
rect 1158 439 1207 753
rect 1534 701 1571 753
rect 1620 800 1669 1471
rect 1791 976 1802 1606
rect 1878 1606 2463 1657
rect 1878 976 1888 1606
rect 1791 964 1888 976
rect 2009 919 2080 1039
rect 2009 861 2080 867
rect 1620 751 1792 800
rect 1490 664 1680 701
rect 1490 500 1527 664
rect 1643 500 1680 664
rect 1201 -45 1207 439
rect 1158 -57 1207 -45
rect 1375 440 1448 451
rect 1375 -44 1382 440
rect 1436 -44 1448 440
rect 1375 -61 1448 -44
rect 1552 -92 1624 451
rect 1743 440 1792 751
rect 1786 -44 1792 440
rect 1743 -59 1792 -44
rect 326 -185 2478 -92
rect 326 -358 537 -185
rect 2337 -358 2478 -185
rect 326 -368 2478 -358
rect 904 -449 959 -397
rect 1040 -449 1046 -397
rect 904 -453 1046 -449
rect 745 -1042 867 -1036
rect 745 -1197 751 -1042
rect 333 -1395 751 -1197
rect 860 -1395 867 -1042
rect 333 -1397 867 -1395
rect 745 -1405 867 -1397
rect 904 -1667 939 -453
rect 1370 -455 1376 -402
rect 1457 -455 1525 -402
rect 1370 -458 1525 -455
rect 1190 -501 1292 -495
rect 1190 -885 1196 -501
rect 1286 -885 1292 -501
rect 1190 -891 1292 -885
rect 977 -1041 1099 -1035
rect 977 -1394 984 -1041
rect 1093 -1394 1099 -1041
rect 977 -1400 1099 -1394
rect 1350 -1414 1356 -1048
rect 1446 -1414 1452 -1048
rect 1489 -1549 1525 -458
rect 1562 -501 1664 -495
rect 1562 -885 1568 -501
rect 1658 -885 1664 -501
rect 1755 -511 1876 -505
rect 1755 -864 1761 -511
rect 1870 -864 1876 -511
rect 1755 -870 1876 -864
rect 1988 -511 2109 -505
rect 1988 -864 1994 -511
rect 2103 -864 2109 -511
rect 1988 -870 2109 -864
rect 1562 -891 1664 -885
rect 2209 -1396 2526 -1196
rect 2209 -1402 2393 -1396
rect 1334 -1579 1685 -1549
rect 1334 -1585 1623 -1579
rect 1617 -1639 1623 -1585
rect 1679 -1639 1685 -1579
rect 1913 -1667 1948 -1460
rect 904 -1715 1948 -1667
rect 1051 -1845 1128 -1837
rect 1051 -1907 1128 -1901
rect 1051 -2061 1087 -1907
rect 894 -2089 1087 -2061
rect 1479 -2064 1515 -1715
rect 1728 -1845 1805 -1839
rect 1728 -1909 1805 -1901
rect 887 -2097 1087 -2089
rect 740 -2148 856 -2142
rect 740 -2285 746 -2148
rect 850 -2285 856 -2148
rect 740 -2291 856 -2285
rect 887 -2584 923 -2097
rect 1322 -2100 1515 -2064
rect 1756 -2062 1792 -1909
rect 2209 -2026 2217 -1402
rect 2387 -2026 2393 -1402
rect 2209 -2036 2393 -2026
rect 1756 -2098 1949 -2062
rect 967 -2148 1083 -2142
rect 967 -2285 973 -2148
rect 1077 -2285 1083 -2148
rect 967 -2291 1083 -2285
rect 1323 -2158 1440 -2152
rect 1323 -2282 1329 -2158
rect 1434 -2282 1440 -2158
rect 1323 -2288 1440 -2282
rect 1166 -2387 1282 -2381
rect 1166 -2524 1172 -2387
rect 1276 -2524 1282 -2387
rect 1166 -2530 1282 -2524
rect 1479 -2573 1515 -2100
rect 1552 -2387 1668 -2381
rect 1552 -2524 1558 -2387
rect 1662 -2524 1668 -2387
rect 1552 -2530 1668 -2524
rect 1750 -2387 1866 -2381
rect 1750 -2524 1756 -2387
rect 1860 -2524 1866 -2387
rect 1750 -2530 1866 -2524
rect 1347 -2609 1515 -2573
rect 1910 -2586 1946 -2098
rect 1978 -2387 2094 -2381
rect 1978 -2524 1984 -2387
rect 2088 -2524 2094 -2387
rect 1978 -2530 2094 -2524
rect 328 -2679 2515 -2670
rect 328 -2898 542 -2679
rect 840 -2711 2515 -2679
rect 2327 -2881 2515 -2711
rect 840 -2898 2515 -2881
rect 328 -2905 2515 -2898
<< via1 >>
rect 544 1622 842 1841
rect 894 867 972 919
rect 803 -46 857 438
rect 2009 867 2080 919
rect 1147 -45 1201 439
rect 1382 -44 1436 440
rect 1732 -44 1786 440
rect 959 -449 1040 -397
rect 751 -1395 860 -1042
rect 1376 -455 1457 -402
rect 1196 -885 1286 -501
rect 984 -1394 1093 -1041
rect 1356 -1414 1446 -1048
rect 1568 -885 1658 -501
rect 1761 -864 1870 -511
rect 1994 -864 2103 -511
rect 1623 -1639 1679 -1579
rect 1051 -1901 1128 -1845
rect 1728 -1901 1805 -1845
rect 746 -2285 850 -2148
rect 2217 -2026 2387 -1402
rect 973 -2285 1077 -2148
rect 1329 -2282 1434 -2158
rect 1172 -2524 1276 -2387
rect 1558 -2524 1662 -2387
rect 1756 -2524 1860 -2387
rect 1984 -2524 2088 -2387
rect 542 -2711 840 -2679
rect 542 -2881 582 -2711
rect 582 -2881 840 -2711
rect 542 -2898 840 -2881
<< metal2 >>
rect 529 1841 867 1856
rect 529 1622 544 1841
rect 842 1622 867 1841
rect 529 1606 867 1622
rect 529 -2670 660 1606
rect 886 867 894 919
rect 972 867 2009 919
rect 2080 867 2087 919
rect 795 439 1207 441
rect 795 438 1147 439
rect 795 -46 803 438
rect 857 -45 1147 438
rect 1201 -45 1207 439
rect 857 -46 1207 -45
rect 795 -47 1207 -46
rect 1376 440 1792 442
rect 1376 -44 1382 440
rect 1436 -44 1732 440
rect 1786 -44 1792 440
rect 1376 -46 1792 -44
rect 959 -397 1040 -47
rect 959 -455 1040 -449
rect 1376 -402 1457 -46
rect 1376 -461 1457 -455
rect 736 -501 2393 -489
rect 736 -885 1196 -501
rect 1286 -885 1568 -501
rect 1658 -511 2393 -501
rect 1658 -864 1761 -511
rect 1870 -864 1994 -511
rect 2103 -864 2393 -511
rect 1658 -885 2393 -864
rect 736 -893 2393 -885
rect 732 -1041 2127 -1034
rect 732 -1042 984 -1041
rect 732 -1395 751 -1042
rect 860 -1394 984 -1042
rect 1093 -1048 2127 -1041
rect 1093 -1394 1356 -1048
rect 860 -1395 1356 -1394
rect 732 -1414 1356 -1395
rect 1446 -1414 2127 -1048
rect 2208 -1213 2393 -893
rect 732 -1438 2127 -1414
rect 2209 -1402 2393 -1213
rect 732 -2113 891 -1438
rect 1623 -1579 1679 -1572
rect 1623 -1845 1679 -1639
rect 1043 -1901 1051 -1845
rect 1128 -1901 1728 -1845
rect 1805 -1901 1816 -1845
rect 2209 -2026 2217 -1402
rect 2387 -2026 2393 -1402
rect 732 -2148 2122 -2113
rect 732 -2285 746 -2148
rect 850 -2285 973 -2148
rect 1077 -2158 2122 -2148
rect 1077 -2282 1329 -2158
rect 1434 -2282 2122 -2158
rect 1077 -2285 2122 -2282
rect 732 -2297 2122 -2285
rect 2209 -2358 2393 -2026
rect 733 -2387 2393 -2358
rect 733 -2524 1172 -2387
rect 1276 -2524 1558 -2387
rect 1662 -2524 1756 -2387
rect 1860 -2524 1984 -2387
rect 2088 -2524 2393 -2387
rect 733 -2542 2393 -2524
rect 529 -2679 849 -2670
rect 529 -2898 542 -2679
rect 840 -2898 849 -2679
rect 529 -2905 849 -2898
use sky130_fd_pr__pfet_g5v0d10v5_GTJ6Y6  sky130_fd_pr__pfet_g5v0d10v5_GTJ6Y6_0 paramcells
timestamp 1718242007
transform 1 0 1585 0 -1 232
box -387 -512 387 512
use sky130_fd_pr__pfet_g5v0d10v5_U6NWY6  sky130_fd_pr__pfet_g5v0d10v5_U6NWY6_0 paramcells
timestamp 1718242347
transform 1 0 1427 0 1 -1038
box -387 -762 387 762
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  sky130_fd_pr__pfet_g5v0d10v5_U62SY6_0 paramcells
timestamp 1718242097
transform 1 0 1932 0 1 -1038
box -308 -762 308 762
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  sky130_fd_pr__pfet_g5v0d10v5_U62SY6_1
timestamp 1718242097
transform 1 0 922 0 1 -1038
box -308 -762 308 762
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XD1 paramcells
timestamp 1718245724
transform 1 0 2045 0 -1 1003
box -183 -183 183 183
use sky130_fd_pr__nfet_g5v0d10v5_EJGQFX  XM1 paramcells
timestamp 1718245724
transform -1 0 1417 0 1 -2336
box -357 -458 357 458
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM3 paramcells
timestamp 1718245724
transform -1 0 907 0 1 -2336
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM5
timestamp 1718245724
transform 1 0 1927 0 1 -2336
box -278 -458 278 458
use sky130_fd_pr__pfet_g5v0d10v5_GTJ6Y6  XM7
timestamp 1718242007
transform 1 0 1001 0 -1 232
box -387 -512 387 512
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM8
timestamp 1718245724
transform 1 0 964 0 -1 1266
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM10
timestamp 1718245724
transform 1 0 1546 0 -1 1266
box -278 -458 278 458
<< labels >>
flabel metal1 326 -352 526 -152 0 FreeSans 256 0 0 0 vdd
port 5 nsew
flabel metal1 1705 773 1705 773 0 FreeSans 320 0 0 0 holdp
flabel metal1 1271 778 1271 778 0 FreeSans 320 0 0 0 holdb
flabel metal1 340 790 540 990 0 FreeSans 256 0 0 0 hold
port 1 nsew
flabel metal1 336 -2891 536 -2691 0 FreeSans 256 0 0 0 vss
port 2 nsew
flabel metal1 2326 -1396 2526 -1196 0 FreeSans 256 0 0 0 out
port 3 nsew
flabel metal1 333 -1397 533 -1197 0 FreeSans 256 0 0 0 in
port 4 nsew
<< end >>
