magic
tech sky130A
magscale 1 2
timestamp 1717690002
<< nwell >>
rect -4653 -1269 4653 1269
<< mvpmos >>
rect -4395 772 -4295 972
rect -4237 772 -4137 972
rect -4079 772 -3979 972
rect -3921 772 -3821 972
rect -3763 772 -3663 972
rect -3605 772 -3505 972
rect -3447 772 -3347 972
rect -3289 772 -3189 972
rect -3131 772 -3031 972
rect -2973 772 -2873 972
rect -2815 772 -2715 972
rect -2657 772 -2557 972
rect -2499 772 -2399 972
rect -2341 772 -2241 972
rect -2183 772 -2083 972
rect -2025 772 -1925 972
rect -1867 772 -1767 972
rect -1709 772 -1609 972
rect -1551 772 -1451 972
rect -1393 772 -1293 972
rect -1235 772 -1135 972
rect -1077 772 -977 972
rect -919 772 -819 972
rect -761 772 -661 972
rect -603 772 -503 972
rect -445 772 -345 972
rect -287 772 -187 972
rect -129 772 -29 972
rect 29 772 129 972
rect 187 772 287 972
rect 345 772 445 972
rect 503 772 603 972
rect 661 772 761 972
rect 819 772 919 972
rect 977 772 1077 972
rect 1135 772 1235 972
rect 1293 772 1393 972
rect 1451 772 1551 972
rect 1609 772 1709 972
rect 1767 772 1867 972
rect 1925 772 2025 972
rect 2083 772 2183 972
rect 2241 772 2341 972
rect 2399 772 2499 972
rect 2557 772 2657 972
rect 2715 772 2815 972
rect 2873 772 2973 972
rect 3031 772 3131 972
rect 3189 772 3289 972
rect 3347 772 3447 972
rect 3505 772 3605 972
rect 3663 772 3763 972
rect 3821 772 3921 972
rect 3979 772 4079 972
rect 4137 772 4237 972
rect 4295 772 4395 972
rect -4395 336 -4295 536
rect -4237 336 -4137 536
rect -4079 336 -3979 536
rect -3921 336 -3821 536
rect -3763 336 -3663 536
rect -3605 336 -3505 536
rect -3447 336 -3347 536
rect -3289 336 -3189 536
rect -3131 336 -3031 536
rect -2973 336 -2873 536
rect -2815 336 -2715 536
rect -2657 336 -2557 536
rect -2499 336 -2399 536
rect -2341 336 -2241 536
rect -2183 336 -2083 536
rect -2025 336 -1925 536
rect -1867 336 -1767 536
rect -1709 336 -1609 536
rect -1551 336 -1451 536
rect -1393 336 -1293 536
rect -1235 336 -1135 536
rect -1077 336 -977 536
rect -919 336 -819 536
rect -761 336 -661 536
rect -603 336 -503 536
rect -445 336 -345 536
rect -287 336 -187 536
rect -129 336 -29 536
rect 29 336 129 536
rect 187 336 287 536
rect 345 336 445 536
rect 503 336 603 536
rect 661 336 761 536
rect 819 336 919 536
rect 977 336 1077 536
rect 1135 336 1235 536
rect 1293 336 1393 536
rect 1451 336 1551 536
rect 1609 336 1709 536
rect 1767 336 1867 536
rect 1925 336 2025 536
rect 2083 336 2183 536
rect 2241 336 2341 536
rect 2399 336 2499 536
rect 2557 336 2657 536
rect 2715 336 2815 536
rect 2873 336 2973 536
rect 3031 336 3131 536
rect 3189 336 3289 536
rect 3347 336 3447 536
rect 3505 336 3605 536
rect 3663 336 3763 536
rect 3821 336 3921 536
rect 3979 336 4079 536
rect 4137 336 4237 536
rect 4295 336 4395 536
rect -4395 -100 -4295 100
rect -4237 -100 -4137 100
rect -4079 -100 -3979 100
rect -3921 -100 -3821 100
rect -3763 -100 -3663 100
rect -3605 -100 -3505 100
rect -3447 -100 -3347 100
rect -3289 -100 -3189 100
rect -3131 -100 -3031 100
rect -2973 -100 -2873 100
rect -2815 -100 -2715 100
rect -2657 -100 -2557 100
rect -2499 -100 -2399 100
rect -2341 -100 -2241 100
rect -2183 -100 -2083 100
rect -2025 -100 -1925 100
rect -1867 -100 -1767 100
rect -1709 -100 -1609 100
rect -1551 -100 -1451 100
rect -1393 -100 -1293 100
rect -1235 -100 -1135 100
rect -1077 -100 -977 100
rect -919 -100 -819 100
rect -761 -100 -661 100
rect -603 -100 -503 100
rect -445 -100 -345 100
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
rect 345 -100 445 100
rect 503 -100 603 100
rect 661 -100 761 100
rect 819 -100 919 100
rect 977 -100 1077 100
rect 1135 -100 1235 100
rect 1293 -100 1393 100
rect 1451 -100 1551 100
rect 1609 -100 1709 100
rect 1767 -100 1867 100
rect 1925 -100 2025 100
rect 2083 -100 2183 100
rect 2241 -100 2341 100
rect 2399 -100 2499 100
rect 2557 -100 2657 100
rect 2715 -100 2815 100
rect 2873 -100 2973 100
rect 3031 -100 3131 100
rect 3189 -100 3289 100
rect 3347 -100 3447 100
rect 3505 -100 3605 100
rect 3663 -100 3763 100
rect 3821 -100 3921 100
rect 3979 -100 4079 100
rect 4137 -100 4237 100
rect 4295 -100 4395 100
rect -4395 -536 -4295 -336
rect -4237 -536 -4137 -336
rect -4079 -536 -3979 -336
rect -3921 -536 -3821 -336
rect -3763 -536 -3663 -336
rect -3605 -536 -3505 -336
rect -3447 -536 -3347 -336
rect -3289 -536 -3189 -336
rect -3131 -536 -3031 -336
rect -2973 -536 -2873 -336
rect -2815 -536 -2715 -336
rect -2657 -536 -2557 -336
rect -2499 -536 -2399 -336
rect -2341 -536 -2241 -336
rect -2183 -536 -2083 -336
rect -2025 -536 -1925 -336
rect -1867 -536 -1767 -336
rect -1709 -536 -1609 -336
rect -1551 -536 -1451 -336
rect -1393 -536 -1293 -336
rect -1235 -536 -1135 -336
rect -1077 -536 -977 -336
rect -919 -536 -819 -336
rect -761 -536 -661 -336
rect -603 -536 -503 -336
rect -445 -536 -345 -336
rect -287 -536 -187 -336
rect -129 -536 -29 -336
rect 29 -536 129 -336
rect 187 -536 287 -336
rect 345 -536 445 -336
rect 503 -536 603 -336
rect 661 -536 761 -336
rect 819 -536 919 -336
rect 977 -536 1077 -336
rect 1135 -536 1235 -336
rect 1293 -536 1393 -336
rect 1451 -536 1551 -336
rect 1609 -536 1709 -336
rect 1767 -536 1867 -336
rect 1925 -536 2025 -336
rect 2083 -536 2183 -336
rect 2241 -536 2341 -336
rect 2399 -536 2499 -336
rect 2557 -536 2657 -336
rect 2715 -536 2815 -336
rect 2873 -536 2973 -336
rect 3031 -536 3131 -336
rect 3189 -536 3289 -336
rect 3347 -536 3447 -336
rect 3505 -536 3605 -336
rect 3663 -536 3763 -336
rect 3821 -536 3921 -336
rect 3979 -536 4079 -336
rect 4137 -536 4237 -336
rect 4295 -536 4395 -336
rect -4395 -972 -4295 -772
rect -4237 -972 -4137 -772
rect -4079 -972 -3979 -772
rect -3921 -972 -3821 -772
rect -3763 -972 -3663 -772
rect -3605 -972 -3505 -772
rect -3447 -972 -3347 -772
rect -3289 -972 -3189 -772
rect -3131 -972 -3031 -772
rect -2973 -972 -2873 -772
rect -2815 -972 -2715 -772
rect -2657 -972 -2557 -772
rect -2499 -972 -2399 -772
rect -2341 -972 -2241 -772
rect -2183 -972 -2083 -772
rect -2025 -972 -1925 -772
rect -1867 -972 -1767 -772
rect -1709 -972 -1609 -772
rect -1551 -972 -1451 -772
rect -1393 -972 -1293 -772
rect -1235 -972 -1135 -772
rect -1077 -972 -977 -772
rect -919 -972 -819 -772
rect -761 -972 -661 -772
rect -603 -972 -503 -772
rect -445 -972 -345 -772
rect -287 -972 -187 -772
rect -129 -972 -29 -772
rect 29 -972 129 -772
rect 187 -972 287 -772
rect 345 -972 445 -772
rect 503 -972 603 -772
rect 661 -972 761 -772
rect 819 -972 919 -772
rect 977 -972 1077 -772
rect 1135 -972 1235 -772
rect 1293 -972 1393 -772
rect 1451 -972 1551 -772
rect 1609 -972 1709 -772
rect 1767 -972 1867 -772
rect 1925 -972 2025 -772
rect 2083 -972 2183 -772
rect 2241 -972 2341 -772
rect 2399 -972 2499 -772
rect 2557 -972 2657 -772
rect 2715 -972 2815 -772
rect 2873 -972 2973 -772
rect 3031 -972 3131 -772
rect 3189 -972 3289 -772
rect 3347 -972 3447 -772
rect 3505 -972 3605 -772
rect 3663 -972 3763 -772
rect 3821 -972 3921 -772
rect 3979 -972 4079 -772
rect 4137 -972 4237 -772
rect 4295 -972 4395 -772
<< mvpdiff >>
rect -4453 960 -4395 972
rect -4453 784 -4441 960
rect -4407 784 -4395 960
rect -4453 772 -4395 784
rect -4295 960 -4237 972
rect -4295 784 -4283 960
rect -4249 784 -4237 960
rect -4295 772 -4237 784
rect -4137 960 -4079 972
rect -4137 784 -4125 960
rect -4091 784 -4079 960
rect -4137 772 -4079 784
rect -3979 960 -3921 972
rect -3979 784 -3967 960
rect -3933 784 -3921 960
rect -3979 772 -3921 784
rect -3821 960 -3763 972
rect -3821 784 -3809 960
rect -3775 784 -3763 960
rect -3821 772 -3763 784
rect -3663 960 -3605 972
rect -3663 784 -3651 960
rect -3617 784 -3605 960
rect -3663 772 -3605 784
rect -3505 960 -3447 972
rect -3505 784 -3493 960
rect -3459 784 -3447 960
rect -3505 772 -3447 784
rect -3347 960 -3289 972
rect -3347 784 -3335 960
rect -3301 784 -3289 960
rect -3347 772 -3289 784
rect -3189 960 -3131 972
rect -3189 784 -3177 960
rect -3143 784 -3131 960
rect -3189 772 -3131 784
rect -3031 960 -2973 972
rect -3031 784 -3019 960
rect -2985 784 -2973 960
rect -3031 772 -2973 784
rect -2873 960 -2815 972
rect -2873 784 -2861 960
rect -2827 784 -2815 960
rect -2873 772 -2815 784
rect -2715 960 -2657 972
rect -2715 784 -2703 960
rect -2669 784 -2657 960
rect -2715 772 -2657 784
rect -2557 960 -2499 972
rect -2557 784 -2545 960
rect -2511 784 -2499 960
rect -2557 772 -2499 784
rect -2399 960 -2341 972
rect -2399 784 -2387 960
rect -2353 784 -2341 960
rect -2399 772 -2341 784
rect -2241 960 -2183 972
rect -2241 784 -2229 960
rect -2195 784 -2183 960
rect -2241 772 -2183 784
rect -2083 960 -2025 972
rect -2083 784 -2071 960
rect -2037 784 -2025 960
rect -2083 772 -2025 784
rect -1925 960 -1867 972
rect -1925 784 -1913 960
rect -1879 784 -1867 960
rect -1925 772 -1867 784
rect -1767 960 -1709 972
rect -1767 784 -1755 960
rect -1721 784 -1709 960
rect -1767 772 -1709 784
rect -1609 960 -1551 972
rect -1609 784 -1597 960
rect -1563 784 -1551 960
rect -1609 772 -1551 784
rect -1451 960 -1393 972
rect -1451 784 -1439 960
rect -1405 784 -1393 960
rect -1451 772 -1393 784
rect -1293 960 -1235 972
rect -1293 784 -1281 960
rect -1247 784 -1235 960
rect -1293 772 -1235 784
rect -1135 960 -1077 972
rect -1135 784 -1123 960
rect -1089 784 -1077 960
rect -1135 772 -1077 784
rect -977 960 -919 972
rect -977 784 -965 960
rect -931 784 -919 960
rect -977 772 -919 784
rect -819 960 -761 972
rect -819 784 -807 960
rect -773 784 -761 960
rect -819 772 -761 784
rect -661 960 -603 972
rect -661 784 -649 960
rect -615 784 -603 960
rect -661 772 -603 784
rect -503 960 -445 972
rect -503 784 -491 960
rect -457 784 -445 960
rect -503 772 -445 784
rect -345 960 -287 972
rect -345 784 -333 960
rect -299 784 -287 960
rect -345 772 -287 784
rect -187 960 -129 972
rect -187 784 -175 960
rect -141 784 -129 960
rect -187 772 -129 784
rect -29 960 29 972
rect -29 784 -17 960
rect 17 784 29 960
rect -29 772 29 784
rect 129 960 187 972
rect 129 784 141 960
rect 175 784 187 960
rect 129 772 187 784
rect 287 960 345 972
rect 287 784 299 960
rect 333 784 345 960
rect 287 772 345 784
rect 445 960 503 972
rect 445 784 457 960
rect 491 784 503 960
rect 445 772 503 784
rect 603 960 661 972
rect 603 784 615 960
rect 649 784 661 960
rect 603 772 661 784
rect 761 960 819 972
rect 761 784 773 960
rect 807 784 819 960
rect 761 772 819 784
rect 919 960 977 972
rect 919 784 931 960
rect 965 784 977 960
rect 919 772 977 784
rect 1077 960 1135 972
rect 1077 784 1089 960
rect 1123 784 1135 960
rect 1077 772 1135 784
rect 1235 960 1293 972
rect 1235 784 1247 960
rect 1281 784 1293 960
rect 1235 772 1293 784
rect 1393 960 1451 972
rect 1393 784 1405 960
rect 1439 784 1451 960
rect 1393 772 1451 784
rect 1551 960 1609 972
rect 1551 784 1563 960
rect 1597 784 1609 960
rect 1551 772 1609 784
rect 1709 960 1767 972
rect 1709 784 1721 960
rect 1755 784 1767 960
rect 1709 772 1767 784
rect 1867 960 1925 972
rect 1867 784 1879 960
rect 1913 784 1925 960
rect 1867 772 1925 784
rect 2025 960 2083 972
rect 2025 784 2037 960
rect 2071 784 2083 960
rect 2025 772 2083 784
rect 2183 960 2241 972
rect 2183 784 2195 960
rect 2229 784 2241 960
rect 2183 772 2241 784
rect 2341 960 2399 972
rect 2341 784 2353 960
rect 2387 784 2399 960
rect 2341 772 2399 784
rect 2499 960 2557 972
rect 2499 784 2511 960
rect 2545 784 2557 960
rect 2499 772 2557 784
rect 2657 960 2715 972
rect 2657 784 2669 960
rect 2703 784 2715 960
rect 2657 772 2715 784
rect 2815 960 2873 972
rect 2815 784 2827 960
rect 2861 784 2873 960
rect 2815 772 2873 784
rect 2973 960 3031 972
rect 2973 784 2985 960
rect 3019 784 3031 960
rect 2973 772 3031 784
rect 3131 960 3189 972
rect 3131 784 3143 960
rect 3177 784 3189 960
rect 3131 772 3189 784
rect 3289 960 3347 972
rect 3289 784 3301 960
rect 3335 784 3347 960
rect 3289 772 3347 784
rect 3447 960 3505 972
rect 3447 784 3459 960
rect 3493 784 3505 960
rect 3447 772 3505 784
rect 3605 960 3663 972
rect 3605 784 3617 960
rect 3651 784 3663 960
rect 3605 772 3663 784
rect 3763 960 3821 972
rect 3763 784 3775 960
rect 3809 784 3821 960
rect 3763 772 3821 784
rect 3921 960 3979 972
rect 3921 784 3933 960
rect 3967 784 3979 960
rect 3921 772 3979 784
rect 4079 960 4137 972
rect 4079 784 4091 960
rect 4125 784 4137 960
rect 4079 772 4137 784
rect 4237 960 4295 972
rect 4237 784 4249 960
rect 4283 784 4295 960
rect 4237 772 4295 784
rect 4395 960 4453 972
rect 4395 784 4407 960
rect 4441 784 4453 960
rect 4395 772 4453 784
rect -4453 524 -4395 536
rect -4453 348 -4441 524
rect -4407 348 -4395 524
rect -4453 336 -4395 348
rect -4295 524 -4237 536
rect -4295 348 -4283 524
rect -4249 348 -4237 524
rect -4295 336 -4237 348
rect -4137 524 -4079 536
rect -4137 348 -4125 524
rect -4091 348 -4079 524
rect -4137 336 -4079 348
rect -3979 524 -3921 536
rect -3979 348 -3967 524
rect -3933 348 -3921 524
rect -3979 336 -3921 348
rect -3821 524 -3763 536
rect -3821 348 -3809 524
rect -3775 348 -3763 524
rect -3821 336 -3763 348
rect -3663 524 -3605 536
rect -3663 348 -3651 524
rect -3617 348 -3605 524
rect -3663 336 -3605 348
rect -3505 524 -3447 536
rect -3505 348 -3493 524
rect -3459 348 -3447 524
rect -3505 336 -3447 348
rect -3347 524 -3289 536
rect -3347 348 -3335 524
rect -3301 348 -3289 524
rect -3347 336 -3289 348
rect -3189 524 -3131 536
rect -3189 348 -3177 524
rect -3143 348 -3131 524
rect -3189 336 -3131 348
rect -3031 524 -2973 536
rect -3031 348 -3019 524
rect -2985 348 -2973 524
rect -3031 336 -2973 348
rect -2873 524 -2815 536
rect -2873 348 -2861 524
rect -2827 348 -2815 524
rect -2873 336 -2815 348
rect -2715 524 -2657 536
rect -2715 348 -2703 524
rect -2669 348 -2657 524
rect -2715 336 -2657 348
rect -2557 524 -2499 536
rect -2557 348 -2545 524
rect -2511 348 -2499 524
rect -2557 336 -2499 348
rect -2399 524 -2341 536
rect -2399 348 -2387 524
rect -2353 348 -2341 524
rect -2399 336 -2341 348
rect -2241 524 -2183 536
rect -2241 348 -2229 524
rect -2195 348 -2183 524
rect -2241 336 -2183 348
rect -2083 524 -2025 536
rect -2083 348 -2071 524
rect -2037 348 -2025 524
rect -2083 336 -2025 348
rect -1925 524 -1867 536
rect -1925 348 -1913 524
rect -1879 348 -1867 524
rect -1925 336 -1867 348
rect -1767 524 -1709 536
rect -1767 348 -1755 524
rect -1721 348 -1709 524
rect -1767 336 -1709 348
rect -1609 524 -1551 536
rect -1609 348 -1597 524
rect -1563 348 -1551 524
rect -1609 336 -1551 348
rect -1451 524 -1393 536
rect -1451 348 -1439 524
rect -1405 348 -1393 524
rect -1451 336 -1393 348
rect -1293 524 -1235 536
rect -1293 348 -1281 524
rect -1247 348 -1235 524
rect -1293 336 -1235 348
rect -1135 524 -1077 536
rect -1135 348 -1123 524
rect -1089 348 -1077 524
rect -1135 336 -1077 348
rect -977 524 -919 536
rect -977 348 -965 524
rect -931 348 -919 524
rect -977 336 -919 348
rect -819 524 -761 536
rect -819 348 -807 524
rect -773 348 -761 524
rect -819 336 -761 348
rect -661 524 -603 536
rect -661 348 -649 524
rect -615 348 -603 524
rect -661 336 -603 348
rect -503 524 -445 536
rect -503 348 -491 524
rect -457 348 -445 524
rect -503 336 -445 348
rect -345 524 -287 536
rect -345 348 -333 524
rect -299 348 -287 524
rect -345 336 -287 348
rect -187 524 -129 536
rect -187 348 -175 524
rect -141 348 -129 524
rect -187 336 -129 348
rect -29 524 29 536
rect -29 348 -17 524
rect 17 348 29 524
rect -29 336 29 348
rect 129 524 187 536
rect 129 348 141 524
rect 175 348 187 524
rect 129 336 187 348
rect 287 524 345 536
rect 287 348 299 524
rect 333 348 345 524
rect 287 336 345 348
rect 445 524 503 536
rect 445 348 457 524
rect 491 348 503 524
rect 445 336 503 348
rect 603 524 661 536
rect 603 348 615 524
rect 649 348 661 524
rect 603 336 661 348
rect 761 524 819 536
rect 761 348 773 524
rect 807 348 819 524
rect 761 336 819 348
rect 919 524 977 536
rect 919 348 931 524
rect 965 348 977 524
rect 919 336 977 348
rect 1077 524 1135 536
rect 1077 348 1089 524
rect 1123 348 1135 524
rect 1077 336 1135 348
rect 1235 524 1293 536
rect 1235 348 1247 524
rect 1281 348 1293 524
rect 1235 336 1293 348
rect 1393 524 1451 536
rect 1393 348 1405 524
rect 1439 348 1451 524
rect 1393 336 1451 348
rect 1551 524 1609 536
rect 1551 348 1563 524
rect 1597 348 1609 524
rect 1551 336 1609 348
rect 1709 524 1767 536
rect 1709 348 1721 524
rect 1755 348 1767 524
rect 1709 336 1767 348
rect 1867 524 1925 536
rect 1867 348 1879 524
rect 1913 348 1925 524
rect 1867 336 1925 348
rect 2025 524 2083 536
rect 2025 348 2037 524
rect 2071 348 2083 524
rect 2025 336 2083 348
rect 2183 524 2241 536
rect 2183 348 2195 524
rect 2229 348 2241 524
rect 2183 336 2241 348
rect 2341 524 2399 536
rect 2341 348 2353 524
rect 2387 348 2399 524
rect 2341 336 2399 348
rect 2499 524 2557 536
rect 2499 348 2511 524
rect 2545 348 2557 524
rect 2499 336 2557 348
rect 2657 524 2715 536
rect 2657 348 2669 524
rect 2703 348 2715 524
rect 2657 336 2715 348
rect 2815 524 2873 536
rect 2815 348 2827 524
rect 2861 348 2873 524
rect 2815 336 2873 348
rect 2973 524 3031 536
rect 2973 348 2985 524
rect 3019 348 3031 524
rect 2973 336 3031 348
rect 3131 524 3189 536
rect 3131 348 3143 524
rect 3177 348 3189 524
rect 3131 336 3189 348
rect 3289 524 3347 536
rect 3289 348 3301 524
rect 3335 348 3347 524
rect 3289 336 3347 348
rect 3447 524 3505 536
rect 3447 348 3459 524
rect 3493 348 3505 524
rect 3447 336 3505 348
rect 3605 524 3663 536
rect 3605 348 3617 524
rect 3651 348 3663 524
rect 3605 336 3663 348
rect 3763 524 3821 536
rect 3763 348 3775 524
rect 3809 348 3821 524
rect 3763 336 3821 348
rect 3921 524 3979 536
rect 3921 348 3933 524
rect 3967 348 3979 524
rect 3921 336 3979 348
rect 4079 524 4137 536
rect 4079 348 4091 524
rect 4125 348 4137 524
rect 4079 336 4137 348
rect 4237 524 4295 536
rect 4237 348 4249 524
rect 4283 348 4295 524
rect 4237 336 4295 348
rect 4395 524 4453 536
rect 4395 348 4407 524
rect 4441 348 4453 524
rect 4395 336 4453 348
rect -4453 88 -4395 100
rect -4453 -88 -4441 88
rect -4407 -88 -4395 88
rect -4453 -100 -4395 -88
rect -4295 88 -4237 100
rect -4295 -88 -4283 88
rect -4249 -88 -4237 88
rect -4295 -100 -4237 -88
rect -4137 88 -4079 100
rect -4137 -88 -4125 88
rect -4091 -88 -4079 88
rect -4137 -100 -4079 -88
rect -3979 88 -3921 100
rect -3979 -88 -3967 88
rect -3933 -88 -3921 88
rect -3979 -100 -3921 -88
rect -3821 88 -3763 100
rect -3821 -88 -3809 88
rect -3775 -88 -3763 88
rect -3821 -100 -3763 -88
rect -3663 88 -3605 100
rect -3663 -88 -3651 88
rect -3617 -88 -3605 88
rect -3663 -100 -3605 -88
rect -3505 88 -3447 100
rect -3505 -88 -3493 88
rect -3459 -88 -3447 88
rect -3505 -100 -3447 -88
rect -3347 88 -3289 100
rect -3347 -88 -3335 88
rect -3301 -88 -3289 88
rect -3347 -100 -3289 -88
rect -3189 88 -3131 100
rect -3189 -88 -3177 88
rect -3143 -88 -3131 88
rect -3189 -100 -3131 -88
rect -3031 88 -2973 100
rect -3031 -88 -3019 88
rect -2985 -88 -2973 88
rect -3031 -100 -2973 -88
rect -2873 88 -2815 100
rect -2873 -88 -2861 88
rect -2827 -88 -2815 88
rect -2873 -100 -2815 -88
rect -2715 88 -2657 100
rect -2715 -88 -2703 88
rect -2669 -88 -2657 88
rect -2715 -100 -2657 -88
rect -2557 88 -2499 100
rect -2557 -88 -2545 88
rect -2511 -88 -2499 88
rect -2557 -100 -2499 -88
rect -2399 88 -2341 100
rect -2399 -88 -2387 88
rect -2353 -88 -2341 88
rect -2399 -100 -2341 -88
rect -2241 88 -2183 100
rect -2241 -88 -2229 88
rect -2195 -88 -2183 88
rect -2241 -100 -2183 -88
rect -2083 88 -2025 100
rect -2083 -88 -2071 88
rect -2037 -88 -2025 88
rect -2083 -100 -2025 -88
rect -1925 88 -1867 100
rect -1925 -88 -1913 88
rect -1879 -88 -1867 88
rect -1925 -100 -1867 -88
rect -1767 88 -1709 100
rect -1767 -88 -1755 88
rect -1721 -88 -1709 88
rect -1767 -100 -1709 -88
rect -1609 88 -1551 100
rect -1609 -88 -1597 88
rect -1563 -88 -1551 88
rect -1609 -100 -1551 -88
rect -1451 88 -1393 100
rect -1451 -88 -1439 88
rect -1405 -88 -1393 88
rect -1451 -100 -1393 -88
rect -1293 88 -1235 100
rect -1293 -88 -1281 88
rect -1247 -88 -1235 88
rect -1293 -100 -1235 -88
rect -1135 88 -1077 100
rect -1135 -88 -1123 88
rect -1089 -88 -1077 88
rect -1135 -100 -1077 -88
rect -977 88 -919 100
rect -977 -88 -965 88
rect -931 -88 -919 88
rect -977 -100 -919 -88
rect -819 88 -761 100
rect -819 -88 -807 88
rect -773 -88 -761 88
rect -819 -100 -761 -88
rect -661 88 -603 100
rect -661 -88 -649 88
rect -615 -88 -603 88
rect -661 -100 -603 -88
rect -503 88 -445 100
rect -503 -88 -491 88
rect -457 -88 -445 88
rect -503 -100 -445 -88
rect -345 88 -287 100
rect -345 -88 -333 88
rect -299 -88 -287 88
rect -345 -100 -287 -88
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
rect 287 88 345 100
rect 287 -88 299 88
rect 333 -88 345 88
rect 287 -100 345 -88
rect 445 88 503 100
rect 445 -88 457 88
rect 491 -88 503 88
rect 445 -100 503 -88
rect 603 88 661 100
rect 603 -88 615 88
rect 649 -88 661 88
rect 603 -100 661 -88
rect 761 88 819 100
rect 761 -88 773 88
rect 807 -88 819 88
rect 761 -100 819 -88
rect 919 88 977 100
rect 919 -88 931 88
rect 965 -88 977 88
rect 919 -100 977 -88
rect 1077 88 1135 100
rect 1077 -88 1089 88
rect 1123 -88 1135 88
rect 1077 -100 1135 -88
rect 1235 88 1293 100
rect 1235 -88 1247 88
rect 1281 -88 1293 88
rect 1235 -100 1293 -88
rect 1393 88 1451 100
rect 1393 -88 1405 88
rect 1439 -88 1451 88
rect 1393 -100 1451 -88
rect 1551 88 1609 100
rect 1551 -88 1563 88
rect 1597 -88 1609 88
rect 1551 -100 1609 -88
rect 1709 88 1767 100
rect 1709 -88 1721 88
rect 1755 -88 1767 88
rect 1709 -100 1767 -88
rect 1867 88 1925 100
rect 1867 -88 1879 88
rect 1913 -88 1925 88
rect 1867 -100 1925 -88
rect 2025 88 2083 100
rect 2025 -88 2037 88
rect 2071 -88 2083 88
rect 2025 -100 2083 -88
rect 2183 88 2241 100
rect 2183 -88 2195 88
rect 2229 -88 2241 88
rect 2183 -100 2241 -88
rect 2341 88 2399 100
rect 2341 -88 2353 88
rect 2387 -88 2399 88
rect 2341 -100 2399 -88
rect 2499 88 2557 100
rect 2499 -88 2511 88
rect 2545 -88 2557 88
rect 2499 -100 2557 -88
rect 2657 88 2715 100
rect 2657 -88 2669 88
rect 2703 -88 2715 88
rect 2657 -100 2715 -88
rect 2815 88 2873 100
rect 2815 -88 2827 88
rect 2861 -88 2873 88
rect 2815 -100 2873 -88
rect 2973 88 3031 100
rect 2973 -88 2985 88
rect 3019 -88 3031 88
rect 2973 -100 3031 -88
rect 3131 88 3189 100
rect 3131 -88 3143 88
rect 3177 -88 3189 88
rect 3131 -100 3189 -88
rect 3289 88 3347 100
rect 3289 -88 3301 88
rect 3335 -88 3347 88
rect 3289 -100 3347 -88
rect 3447 88 3505 100
rect 3447 -88 3459 88
rect 3493 -88 3505 88
rect 3447 -100 3505 -88
rect 3605 88 3663 100
rect 3605 -88 3617 88
rect 3651 -88 3663 88
rect 3605 -100 3663 -88
rect 3763 88 3821 100
rect 3763 -88 3775 88
rect 3809 -88 3821 88
rect 3763 -100 3821 -88
rect 3921 88 3979 100
rect 3921 -88 3933 88
rect 3967 -88 3979 88
rect 3921 -100 3979 -88
rect 4079 88 4137 100
rect 4079 -88 4091 88
rect 4125 -88 4137 88
rect 4079 -100 4137 -88
rect 4237 88 4295 100
rect 4237 -88 4249 88
rect 4283 -88 4295 88
rect 4237 -100 4295 -88
rect 4395 88 4453 100
rect 4395 -88 4407 88
rect 4441 -88 4453 88
rect 4395 -100 4453 -88
rect -4453 -348 -4395 -336
rect -4453 -524 -4441 -348
rect -4407 -524 -4395 -348
rect -4453 -536 -4395 -524
rect -4295 -348 -4237 -336
rect -4295 -524 -4283 -348
rect -4249 -524 -4237 -348
rect -4295 -536 -4237 -524
rect -4137 -348 -4079 -336
rect -4137 -524 -4125 -348
rect -4091 -524 -4079 -348
rect -4137 -536 -4079 -524
rect -3979 -348 -3921 -336
rect -3979 -524 -3967 -348
rect -3933 -524 -3921 -348
rect -3979 -536 -3921 -524
rect -3821 -348 -3763 -336
rect -3821 -524 -3809 -348
rect -3775 -524 -3763 -348
rect -3821 -536 -3763 -524
rect -3663 -348 -3605 -336
rect -3663 -524 -3651 -348
rect -3617 -524 -3605 -348
rect -3663 -536 -3605 -524
rect -3505 -348 -3447 -336
rect -3505 -524 -3493 -348
rect -3459 -524 -3447 -348
rect -3505 -536 -3447 -524
rect -3347 -348 -3289 -336
rect -3347 -524 -3335 -348
rect -3301 -524 -3289 -348
rect -3347 -536 -3289 -524
rect -3189 -348 -3131 -336
rect -3189 -524 -3177 -348
rect -3143 -524 -3131 -348
rect -3189 -536 -3131 -524
rect -3031 -348 -2973 -336
rect -3031 -524 -3019 -348
rect -2985 -524 -2973 -348
rect -3031 -536 -2973 -524
rect -2873 -348 -2815 -336
rect -2873 -524 -2861 -348
rect -2827 -524 -2815 -348
rect -2873 -536 -2815 -524
rect -2715 -348 -2657 -336
rect -2715 -524 -2703 -348
rect -2669 -524 -2657 -348
rect -2715 -536 -2657 -524
rect -2557 -348 -2499 -336
rect -2557 -524 -2545 -348
rect -2511 -524 -2499 -348
rect -2557 -536 -2499 -524
rect -2399 -348 -2341 -336
rect -2399 -524 -2387 -348
rect -2353 -524 -2341 -348
rect -2399 -536 -2341 -524
rect -2241 -348 -2183 -336
rect -2241 -524 -2229 -348
rect -2195 -524 -2183 -348
rect -2241 -536 -2183 -524
rect -2083 -348 -2025 -336
rect -2083 -524 -2071 -348
rect -2037 -524 -2025 -348
rect -2083 -536 -2025 -524
rect -1925 -348 -1867 -336
rect -1925 -524 -1913 -348
rect -1879 -524 -1867 -348
rect -1925 -536 -1867 -524
rect -1767 -348 -1709 -336
rect -1767 -524 -1755 -348
rect -1721 -524 -1709 -348
rect -1767 -536 -1709 -524
rect -1609 -348 -1551 -336
rect -1609 -524 -1597 -348
rect -1563 -524 -1551 -348
rect -1609 -536 -1551 -524
rect -1451 -348 -1393 -336
rect -1451 -524 -1439 -348
rect -1405 -524 -1393 -348
rect -1451 -536 -1393 -524
rect -1293 -348 -1235 -336
rect -1293 -524 -1281 -348
rect -1247 -524 -1235 -348
rect -1293 -536 -1235 -524
rect -1135 -348 -1077 -336
rect -1135 -524 -1123 -348
rect -1089 -524 -1077 -348
rect -1135 -536 -1077 -524
rect -977 -348 -919 -336
rect -977 -524 -965 -348
rect -931 -524 -919 -348
rect -977 -536 -919 -524
rect -819 -348 -761 -336
rect -819 -524 -807 -348
rect -773 -524 -761 -348
rect -819 -536 -761 -524
rect -661 -348 -603 -336
rect -661 -524 -649 -348
rect -615 -524 -603 -348
rect -661 -536 -603 -524
rect -503 -348 -445 -336
rect -503 -524 -491 -348
rect -457 -524 -445 -348
rect -503 -536 -445 -524
rect -345 -348 -287 -336
rect -345 -524 -333 -348
rect -299 -524 -287 -348
rect -345 -536 -287 -524
rect -187 -348 -129 -336
rect -187 -524 -175 -348
rect -141 -524 -129 -348
rect -187 -536 -129 -524
rect -29 -348 29 -336
rect -29 -524 -17 -348
rect 17 -524 29 -348
rect -29 -536 29 -524
rect 129 -348 187 -336
rect 129 -524 141 -348
rect 175 -524 187 -348
rect 129 -536 187 -524
rect 287 -348 345 -336
rect 287 -524 299 -348
rect 333 -524 345 -348
rect 287 -536 345 -524
rect 445 -348 503 -336
rect 445 -524 457 -348
rect 491 -524 503 -348
rect 445 -536 503 -524
rect 603 -348 661 -336
rect 603 -524 615 -348
rect 649 -524 661 -348
rect 603 -536 661 -524
rect 761 -348 819 -336
rect 761 -524 773 -348
rect 807 -524 819 -348
rect 761 -536 819 -524
rect 919 -348 977 -336
rect 919 -524 931 -348
rect 965 -524 977 -348
rect 919 -536 977 -524
rect 1077 -348 1135 -336
rect 1077 -524 1089 -348
rect 1123 -524 1135 -348
rect 1077 -536 1135 -524
rect 1235 -348 1293 -336
rect 1235 -524 1247 -348
rect 1281 -524 1293 -348
rect 1235 -536 1293 -524
rect 1393 -348 1451 -336
rect 1393 -524 1405 -348
rect 1439 -524 1451 -348
rect 1393 -536 1451 -524
rect 1551 -348 1609 -336
rect 1551 -524 1563 -348
rect 1597 -524 1609 -348
rect 1551 -536 1609 -524
rect 1709 -348 1767 -336
rect 1709 -524 1721 -348
rect 1755 -524 1767 -348
rect 1709 -536 1767 -524
rect 1867 -348 1925 -336
rect 1867 -524 1879 -348
rect 1913 -524 1925 -348
rect 1867 -536 1925 -524
rect 2025 -348 2083 -336
rect 2025 -524 2037 -348
rect 2071 -524 2083 -348
rect 2025 -536 2083 -524
rect 2183 -348 2241 -336
rect 2183 -524 2195 -348
rect 2229 -524 2241 -348
rect 2183 -536 2241 -524
rect 2341 -348 2399 -336
rect 2341 -524 2353 -348
rect 2387 -524 2399 -348
rect 2341 -536 2399 -524
rect 2499 -348 2557 -336
rect 2499 -524 2511 -348
rect 2545 -524 2557 -348
rect 2499 -536 2557 -524
rect 2657 -348 2715 -336
rect 2657 -524 2669 -348
rect 2703 -524 2715 -348
rect 2657 -536 2715 -524
rect 2815 -348 2873 -336
rect 2815 -524 2827 -348
rect 2861 -524 2873 -348
rect 2815 -536 2873 -524
rect 2973 -348 3031 -336
rect 2973 -524 2985 -348
rect 3019 -524 3031 -348
rect 2973 -536 3031 -524
rect 3131 -348 3189 -336
rect 3131 -524 3143 -348
rect 3177 -524 3189 -348
rect 3131 -536 3189 -524
rect 3289 -348 3347 -336
rect 3289 -524 3301 -348
rect 3335 -524 3347 -348
rect 3289 -536 3347 -524
rect 3447 -348 3505 -336
rect 3447 -524 3459 -348
rect 3493 -524 3505 -348
rect 3447 -536 3505 -524
rect 3605 -348 3663 -336
rect 3605 -524 3617 -348
rect 3651 -524 3663 -348
rect 3605 -536 3663 -524
rect 3763 -348 3821 -336
rect 3763 -524 3775 -348
rect 3809 -524 3821 -348
rect 3763 -536 3821 -524
rect 3921 -348 3979 -336
rect 3921 -524 3933 -348
rect 3967 -524 3979 -348
rect 3921 -536 3979 -524
rect 4079 -348 4137 -336
rect 4079 -524 4091 -348
rect 4125 -524 4137 -348
rect 4079 -536 4137 -524
rect 4237 -348 4295 -336
rect 4237 -524 4249 -348
rect 4283 -524 4295 -348
rect 4237 -536 4295 -524
rect 4395 -348 4453 -336
rect 4395 -524 4407 -348
rect 4441 -524 4453 -348
rect 4395 -536 4453 -524
rect -4453 -784 -4395 -772
rect -4453 -960 -4441 -784
rect -4407 -960 -4395 -784
rect -4453 -972 -4395 -960
rect -4295 -784 -4237 -772
rect -4295 -960 -4283 -784
rect -4249 -960 -4237 -784
rect -4295 -972 -4237 -960
rect -4137 -784 -4079 -772
rect -4137 -960 -4125 -784
rect -4091 -960 -4079 -784
rect -4137 -972 -4079 -960
rect -3979 -784 -3921 -772
rect -3979 -960 -3967 -784
rect -3933 -960 -3921 -784
rect -3979 -972 -3921 -960
rect -3821 -784 -3763 -772
rect -3821 -960 -3809 -784
rect -3775 -960 -3763 -784
rect -3821 -972 -3763 -960
rect -3663 -784 -3605 -772
rect -3663 -960 -3651 -784
rect -3617 -960 -3605 -784
rect -3663 -972 -3605 -960
rect -3505 -784 -3447 -772
rect -3505 -960 -3493 -784
rect -3459 -960 -3447 -784
rect -3505 -972 -3447 -960
rect -3347 -784 -3289 -772
rect -3347 -960 -3335 -784
rect -3301 -960 -3289 -784
rect -3347 -972 -3289 -960
rect -3189 -784 -3131 -772
rect -3189 -960 -3177 -784
rect -3143 -960 -3131 -784
rect -3189 -972 -3131 -960
rect -3031 -784 -2973 -772
rect -3031 -960 -3019 -784
rect -2985 -960 -2973 -784
rect -3031 -972 -2973 -960
rect -2873 -784 -2815 -772
rect -2873 -960 -2861 -784
rect -2827 -960 -2815 -784
rect -2873 -972 -2815 -960
rect -2715 -784 -2657 -772
rect -2715 -960 -2703 -784
rect -2669 -960 -2657 -784
rect -2715 -972 -2657 -960
rect -2557 -784 -2499 -772
rect -2557 -960 -2545 -784
rect -2511 -960 -2499 -784
rect -2557 -972 -2499 -960
rect -2399 -784 -2341 -772
rect -2399 -960 -2387 -784
rect -2353 -960 -2341 -784
rect -2399 -972 -2341 -960
rect -2241 -784 -2183 -772
rect -2241 -960 -2229 -784
rect -2195 -960 -2183 -784
rect -2241 -972 -2183 -960
rect -2083 -784 -2025 -772
rect -2083 -960 -2071 -784
rect -2037 -960 -2025 -784
rect -2083 -972 -2025 -960
rect -1925 -784 -1867 -772
rect -1925 -960 -1913 -784
rect -1879 -960 -1867 -784
rect -1925 -972 -1867 -960
rect -1767 -784 -1709 -772
rect -1767 -960 -1755 -784
rect -1721 -960 -1709 -784
rect -1767 -972 -1709 -960
rect -1609 -784 -1551 -772
rect -1609 -960 -1597 -784
rect -1563 -960 -1551 -784
rect -1609 -972 -1551 -960
rect -1451 -784 -1393 -772
rect -1451 -960 -1439 -784
rect -1405 -960 -1393 -784
rect -1451 -972 -1393 -960
rect -1293 -784 -1235 -772
rect -1293 -960 -1281 -784
rect -1247 -960 -1235 -784
rect -1293 -972 -1235 -960
rect -1135 -784 -1077 -772
rect -1135 -960 -1123 -784
rect -1089 -960 -1077 -784
rect -1135 -972 -1077 -960
rect -977 -784 -919 -772
rect -977 -960 -965 -784
rect -931 -960 -919 -784
rect -977 -972 -919 -960
rect -819 -784 -761 -772
rect -819 -960 -807 -784
rect -773 -960 -761 -784
rect -819 -972 -761 -960
rect -661 -784 -603 -772
rect -661 -960 -649 -784
rect -615 -960 -603 -784
rect -661 -972 -603 -960
rect -503 -784 -445 -772
rect -503 -960 -491 -784
rect -457 -960 -445 -784
rect -503 -972 -445 -960
rect -345 -784 -287 -772
rect -345 -960 -333 -784
rect -299 -960 -287 -784
rect -345 -972 -287 -960
rect -187 -784 -129 -772
rect -187 -960 -175 -784
rect -141 -960 -129 -784
rect -187 -972 -129 -960
rect -29 -784 29 -772
rect -29 -960 -17 -784
rect 17 -960 29 -784
rect -29 -972 29 -960
rect 129 -784 187 -772
rect 129 -960 141 -784
rect 175 -960 187 -784
rect 129 -972 187 -960
rect 287 -784 345 -772
rect 287 -960 299 -784
rect 333 -960 345 -784
rect 287 -972 345 -960
rect 445 -784 503 -772
rect 445 -960 457 -784
rect 491 -960 503 -784
rect 445 -972 503 -960
rect 603 -784 661 -772
rect 603 -960 615 -784
rect 649 -960 661 -784
rect 603 -972 661 -960
rect 761 -784 819 -772
rect 761 -960 773 -784
rect 807 -960 819 -784
rect 761 -972 819 -960
rect 919 -784 977 -772
rect 919 -960 931 -784
rect 965 -960 977 -784
rect 919 -972 977 -960
rect 1077 -784 1135 -772
rect 1077 -960 1089 -784
rect 1123 -960 1135 -784
rect 1077 -972 1135 -960
rect 1235 -784 1293 -772
rect 1235 -960 1247 -784
rect 1281 -960 1293 -784
rect 1235 -972 1293 -960
rect 1393 -784 1451 -772
rect 1393 -960 1405 -784
rect 1439 -960 1451 -784
rect 1393 -972 1451 -960
rect 1551 -784 1609 -772
rect 1551 -960 1563 -784
rect 1597 -960 1609 -784
rect 1551 -972 1609 -960
rect 1709 -784 1767 -772
rect 1709 -960 1721 -784
rect 1755 -960 1767 -784
rect 1709 -972 1767 -960
rect 1867 -784 1925 -772
rect 1867 -960 1879 -784
rect 1913 -960 1925 -784
rect 1867 -972 1925 -960
rect 2025 -784 2083 -772
rect 2025 -960 2037 -784
rect 2071 -960 2083 -784
rect 2025 -972 2083 -960
rect 2183 -784 2241 -772
rect 2183 -960 2195 -784
rect 2229 -960 2241 -784
rect 2183 -972 2241 -960
rect 2341 -784 2399 -772
rect 2341 -960 2353 -784
rect 2387 -960 2399 -784
rect 2341 -972 2399 -960
rect 2499 -784 2557 -772
rect 2499 -960 2511 -784
rect 2545 -960 2557 -784
rect 2499 -972 2557 -960
rect 2657 -784 2715 -772
rect 2657 -960 2669 -784
rect 2703 -960 2715 -784
rect 2657 -972 2715 -960
rect 2815 -784 2873 -772
rect 2815 -960 2827 -784
rect 2861 -960 2873 -784
rect 2815 -972 2873 -960
rect 2973 -784 3031 -772
rect 2973 -960 2985 -784
rect 3019 -960 3031 -784
rect 2973 -972 3031 -960
rect 3131 -784 3189 -772
rect 3131 -960 3143 -784
rect 3177 -960 3189 -784
rect 3131 -972 3189 -960
rect 3289 -784 3347 -772
rect 3289 -960 3301 -784
rect 3335 -960 3347 -784
rect 3289 -972 3347 -960
rect 3447 -784 3505 -772
rect 3447 -960 3459 -784
rect 3493 -960 3505 -784
rect 3447 -972 3505 -960
rect 3605 -784 3663 -772
rect 3605 -960 3617 -784
rect 3651 -960 3663 -784
rect 3605 -972 3663 -960
rect 3763 -784 3821 -772
rect 3763 -960 3775 -784
rect 3809 -960 3821 -784
rect 3763 -972 3821 -960
rect 3921 -784 3979 -772
rect 3921 -960 3933 -784
rect 3967 -960 3979 -784
rect 3921 -972 3979 -960
rect 4079 -784 4137 -772
rect 4079 -960 4091 -784
rect 4125 -960 4137 -784
rect 4079 -972 4137 -960
rect 4237 -784 4295 -772
rect 4237 -960 4249 -784
rect 4283 -960 4295 -784
rect 4237 -972 4295 -960
rect 4395 -784 4453 -772
rect 4395 -960 4407 -784
rect 4441 -960 4453 -784
rect 4395 -972 4453 -960
<< mvpdiffc >>
rect -4441 784 -4407 960
rect -4283 784 -4249 960
rect -4125 784 -4091 960
rect -3967 784 -3933 960
rect -3809 784 -3775 960
rect -3651 784 -3617 960
rect -3493 784 -3459 960
rect -3335 784 -3301 960
rect -3177 784 -3143 960
rect -3019 784 -2985 960
rect -2861 784 -2827 960
rect -2703 784 -2669 960
rect -2545 784 -2511 960
rect -2387 784 -2353 960
rect -2229 784 -2195 960
rect -2071 784 -2037 960
rect -1913 784 -1879 960
rect -1755 784 -1721 960
rect -1597 784 -1563 960
rect -1439 784 -1405 960
rect -1281 784 -1247 960
rect -1123 784 -1089 960
rect -965 784 -931 960
rect -807 784 -773 960
rect -649 784 -615 960
rect -491 784 -457 960
rect -333 784 -299 960
rect -175 784 -141 960
rect -17 784 17 960
rect 141 784 175 960
rect 299 784 333 960
rect 457 784 491 960
rect 615 784 649 960
rect 773 784 807 960
rect 931 784 965 960
rect 1089 784 1123 960
rect 1247 784 1281 960
rect 1405 784 1439 960
rect 1563 784 1597 960
rect 1721 784 1755 960
rect 1879 784 1913 960
rect 2037 784 2071 960
rect 2195 784 2229 960
rect 2353 784 2387 960
rect 2511 784 2545 960
rect 2669 784 2703 960
rect 2827 784 2861 960
rect 2985 784 3019 960
rect 3143 784 3177 960
rect 3301 784 3335 960
rect 3459 784 3493 960
rect 3617 784 3651 960
rect 3775 784 3809 960
rect 3933 784 3967 960
rect 4091 784 4125 960
rect 4249 784 4283 960
rect 4407 784 4441 960
rect -4441 348 -4407 524
rect -4283 348 -4249 524
rect -4125 348 -4091 524
rect -3967 348 -3933 524
rect -3809 348 -3775 524
rect -3651 348 -3617 524
rect -3493 348 -3459 524
rect -3335 348 -3301 524
rect -3177 348 -3143 524
rect -3019 348 -2985 524
rect -2861 348 -2827 524
rect -2703 348 -2669 524
rect -2545 348 -2511 524
rect -2387 348 -2353 524
rect -2229 348 -2195 524
rect -2071 348 -2037 524
rect -1913 348 -1879 524
rect -1755 348 -1721 524
rect -1597 348 -1563 524
rect -1439 348 -1405 524
rect -1281 348 -1247 524
rect -1123 348 -1089 524
rect -965 348 -931 524
rect -807 348 -773 524
rect -649 348 -615 524
rect -491 348 -457 524
rect -333 348 -299 524
rect -175 348 -141 524
rect -17 348 17 524
rect 141 348 175 524
rect 299 348 333 524
rect 457 348 491 524
rect 615 348 649 524
rect 773 348 807 524
rect 931 348 965 524
rect 1089 348 1123 524
rect 1247 348 1281 524
rect 1405 348 1439 524
rect 1563 348 1597 524
rect 1721 348 1755 524
rect 1879 348 1913 524
rect 2037 348 2071 524
rect 2195 348 2229 524
rect 2353 348 2387 524
rect 2511 348 2545 524
rect 2669 348 2703 524
rect 2827 348 2861 524
rect 2985 348 3019 524
rect 3143 348 3177 524
rect 3301 348 3335 524
rect 3459 348 3493 524
rect 3617 348 3651 524
rect 3775 348 3809 524
rect 3933 348 3967 524
rect 4091 348 4125 524
rect 4249 348 4283 524
rect 4407 348 4441 524
rect -4441 -88 -4407 88
rect -4283 -88 -4249 88
rect -4125 -88 -4091 88
rect -3967 -88 -3933 88
rect -3809 -88 -3775 88
rect -3651 -88 -3617 88
rect -3493 -88 -3459 88
rect -3335 -88 -3301 88
rect -3177 -88 -3143 88
rect -3019 -88 -2985 88
rect -2861 -88 -2827 88
rect -2703 -88 -2669 88
rect -2545 -88 -2511 88
rect -2387 -88 -2353 88
rect -2229 -88 -2195 88
rect -2071 -88 -2037 88
rect -1913 -88 -1879 88
rect -1755 -88 -1721 88
rect -1597 -88 -1563 88
rect -1439 -88 -1405 88
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
rect 1405 -88 1439 88
rect 1563 -88 1597 88
rect 1721 -88 1755 88
rect 1879 -88 1913 88
rect 2037 -88 2071 88
rect 2195 -88 2229 88
rect 2353 -88 2387 88
rect 2511 -88 2545 88
rect 2669 -88 2703 88
rect 2827 -88 2861 88
rect 2985 -88 3019 88
rect 3143 -88 3177 88
rect 3301 -88 3335 88
rect 3459 -88 3493 88
rect 3617 -88 3651 88
rect 3775 -88 3809 88
rect 3933 -88 3967 88
rect 4091 -88 4125 88
rect 4249 -88 4283 88
rect 4407 -88 4441 88
rect -4441 -524 -4407 -348
rect -4283 -524 -4249 -348
rect -4125 -524 -4091 -348
rect -3967 -524 -3933 -348
rect -3809 -524 -3775 -348
rect -3651 -524 -3617 -348
rect -3493 -524 -3459 -348
rect -3335 -524 -3301 -348
rect -3177 -524 -3143 -348
rect -3019 -524 -2985 -348
rect -2861 -524 -2827 -348
rect -2703 -524 -2669 -348
rect -2545 -524 -2511 -348
rect -2387 -524 -2353 -348
rect -2229 -524 -2195 -348
rect -2071 -524 -2037 -348
rect -1913 -524 -1879 -348
rect -1755 -524 -1721 -348
rect -1597 -524 -1563 -348
rect -1439 -524 -1405 -348
rect -1281 -524 -1247 -348
rect -1123 -524 -1089 -348
rect -965 -524 -931 -348
rect -807 -524 -773 -348
rect -649 -524 -615 -348
rect -491 -524 -457 -348
rect -333 -524 -299 -348
rect -175 -524 -141 -348
rect -17 -524 17 -348
rect 141 -524 175 -348
rect 299 -524 333 -348
rect 457 -524 491 -348
rect 615 -524 649 -348
rect 773 -524 807 -348
rect 931 -524 965 -348
rect 1089 -524 1123 -348
rect 1247 -524 1281 -348
rect 1405 -524 1439 -348
rect 1563 -524 1597 -348
rect 1721 -524 1755 -348
rect 1879 -524 1913 -348
rect 2037 -524 2071 -348
rect 2195 -524 2229 -348
rect 2353 -524 2387 -348
rect 2511 -524 2545 -348
rect 2669 -524 2703 -348
rect 2827 -524 2861 -348
rect 2985 -524 3019 -348
rect 3143 -524 3177 -348
rect 3301 -524 3335 -348
rect 3459 -524 3493 -348
rect 3617 -524 3651 -348
rect 3775 -524 3809 -348
rect 3933 -524 3967 -348
rect 4091 -524 4125 -348
rect 4249 -524 4283 -348
rect 4407 -524 4441 -348
rect -4441 -960 -4407 -784
rect -4283 -960 -4249 -784
rect -4125 -960 -4091 -784
rect -3967 -960 -3933 -784
rect -3809 -960 -3775 -784
rect -3651 -960 -3617 -784
rect -3493 -960 -3459 -784
rect -3335 -960 -3301 -784
rect -3177 -960 -3143 -784
rect -3019 -960 -2985 -784
rect -2861 -960 -2827 -784
rect -2703 -960 -2669 -784
rect -2545 -960 -2511 -784
rect -2387 -960 -2353 -784
rect -2229 -960 -2195 -784
rect -2071 -960 -2037 -784
rect -1913 -960 -1879 -784
rect -1755 -960 -1721 -784
rect -1597 -960 -1563 -784
rect -1439 -960 -1405 -784
rect -1281 -960 -1247 -784
rect -1123 -960 -1089 -784
rect -965 -960 -931 -784
rect -807 -960 -773 -784
rect -649 -960 -615 -784
rect -491 -960 -457 -784
rect -333 -960 -299 -784
rect -175 -960 -141 -784
rect -17 -960 17 -784
rect 141 -960 175 -784
rect 299 -960 333 -784
rect 457 -960 491 -784
rect 615 -960 649 -784
rect 773 -960 807 -784
rect 931 -960 965 -784
rect 1089 -960 1123 -784
rect 1247 -960 1281 -784
rect 1405 -960 1439 -784
rect 1563 -960 1597 -784
rect 1721 -960 1755 -784
rect 1879 -960 1913 -784
rect 2037 -960 2071 -784
rect 2195 -960 2229 -784
rect 2353 -960 2387 -784
rect 2511 -960 2545 -784
rect 2669 -960 2703 -784
rect 2827 -960 2861 -784
rect 2985 -960 3019 -784
rect 3143 -960 3177 -784
rect 3301 -960 3335 -784
rect 3459 -960 3493 -784
rect 3617 -960 3651 -784
rect 3775 -960 3809 -784
rect 3933 -960 3967 -784
rect 4091 -960 4125 -784
rect 4249 -960 4283 -784
rect 4407 -960 4441 -784
<< mvnsubdiff >>
rect -4587 1191 4587 1203
rect -4587 1157 -4479 1191
rect 4479 1157 4587 1191
rect -4587 1145 4587 1157
rect -4587 1095 -4529 1145
rect -4587 -1095 -4575 1095
rect -4541 -1095 -4529 1095
rect 4529 1095 4587 1145
rect -4587 -1145 -4529 -1095
rect 4529 -1095 4541 1095
rect 4575 -1095 4587 1095
rect 4529 -1145 4587 -1095
rect -4587 -1157 4587 -1145
rect -4587 -1191 -4479 -1157
rect 4479 -1191 4587 -1157
rect -4587 -1203 4587 -1191
<< mvnsubdiffcont >>
rect -4479 1157 4479 1191
rect -4575 -1095 -4541 1095
rect 4541 -1095 4575 1095
rect -4479 -1191 4479 -1157
<< poly >>
rect -4395 1053 -4295 1069
rect -4395 1019 -4379 1053
rect -4311 1019 -4295 1053
rect -4395 972 -4295 1019
rect -4237 1053 -4137 1069
rect -4237 1019 -4221 1053
rect -4153 1019 -4137 1053
rect -4237 972 -4137 1019
rect -4079 1053 -3979 1069
rect -4079 1019 -4063 1053
rect -3995 1019 -3979 1053
rect -4079 972 -3979 1019
rect -3921 1053 -3821 1069
rect -3921 1019 -3905 1053
rect -3837 1019 -3821 1053
rect -3921 972 -3821 1019
rect -3763 1053 -3663 1069
rect -3763 1019 -3747 1053
rect -3679 1019 -3663 1053
rect -3763 972 -3663 1019
rect -3605 1053 -3505 1069
rect -3605 1019 -3589 1053
rect -3521 1019 -3505 1053
rect -3605 972 -3505 1019
rect -3447 1053 -3347 1069
rect -3447 1019 -3431 1053
rect -3363 1019 -3347 1053
rect -3447 972 -3347 1019
rect -3289 1053 -3189 1069
rect -3289 1019 -3273 1053
rect -3205 1019 -3189 1053
rect -3289 972 -3189 1019
rect -3131 1053 -3031 1069
rect -3131 1019 -3115 1053
rect -3047 1019 -3031 1053
rect -3131 972 -3031 1019
rect -2973 1053 -2873 1069
rect -2973 1019 -2957 1053
rect -2889 1019 -2873 1053
rect -2973 972 -2873 1019
rect -2815 1053 -2715 1069
rect -2815 1019 -2799 1053
rect -2731 1019 -2715 1053
rect -2815 972 -2715 1019
rect -2657 1053 -2557 1069
rect -2657 1019 -2641 1053
rect -2573 1019 -2557 1053
rect -2657 972 -2557 1019
rect -2499 1053 -2399 1069
rect -2499 1019 -2483 1053
rect -2415 1019 -2399 1053
rect -2499 972 -2399 1019
rect -2341 1053 -2241 1069
rect -2341 1019 -2325 1053
rect -2257 1019 -2241 1053
rect -2341 972 -2241 1019
rect -2183 1053 -2083 1069
rect -2183 1019 -2167 1053
rect -2099 1019 -2083 1053
rect -2183 972 -2083 1019
rect -2025 1053 -1925 1069
rect -2025 1019 -2009 1053
rect -1941 1019 -1925 1053
rect -2025 972 -1925 1019
rect -1867 1053 -1767 1069
rect -1867 1019 -1851 1053
rect -1783 1019 -1767 1053
rect -1867 972 -1767 1019
rect -1709 1053 -1609 1069
rect -1709 1019 -1693 1053
rect -1625 1019 -1609 1053
rect -1709 972 -1609 1019
rect -1551 1053 -1451 1069
rect -1551 1019 -1535 1053
rect -1467 1019 -1451 1053
rect -1551 972 -1451 1019
rect -1393 1053 -1293 1069
rect -1393 1019 -1377 1053
rect -1309 1019 -1293 1053
rect -1393 972 -1293 1019
rect -1235 1053 -1135 1069
rect -1235 1019 -1219 1053
rect -1151 1019 -1135 1053
rect -1235 972 -1135 1019
rect -1077 1053 -977 1069
rect -1077 1019 -1061 1053
rect -993 1019 -977 1053
rect -1077 972 -977 1019
rect -919 1053 -819 1069
rect -919 1019 -903 1053
rect -835 1019 -819 1053
rect -919 972 -819 1019
rect -761 1053 -661 1069
rect -761 1019 -745 1053
rect -677 1019 -661 1053
rect -761 972 -661 1019
rect -603 1053 -503 1069
rect -603 1019 -587 1053
rect -519 1019 -503 1053
rect -603 972 -503 1019
rect -445 1053 -345 1069
rect -445 1019 -429 1053
rect -361 1019 -345 1053
rect -445 972 -345 1019
rect -287 1053 -187 1069
rect -287 1019 -271 1053
rect -203 1019 -187 1053
rect -287 972 -187 1019
rect -129 1053 -29 1069
rect -129 1019 -113 1053
rect -45 1019 -29 1053
rect -129 972 -29 1019
rect 29 1053 129 1069
rect 29 1019 45 1053
rect 113 1019 129 1053
rect 29 972 129 1019
rect 187 1053 287 1069
rect 187 1019 203 1053
rect 271 1019 287 1053
rect 187 972 287 1019
rect 345 1053 445 1069
rect 345 1019 361 1053
rect 429 1019 445 1053
rect 345 972 445 1019
rect 503 1053 603 1069
rect 503 1019 519 1053
rect 587 1019 603 1053
rect 503 972 603 1019
rect 661 1053 761 1069
rect 661 1019 677 1053
rect 745 1019 761 1053
rect 661 972 761 1019
rect 819 1053 919 1069
rect 819 1019 835 1053
rect 903 1019 919 1053
rect 819 972 919 1019
rect 977 1053 1077 1069
rect 977 1019 993 1053
rect 1061 1019 1077 1053
rect 977 972 1077 1019
rect 1135 1053 1235 1069
rect 1135 1019 1151 1053
rect 1219 1019 1235 1053
rect 1135 972 1235 1019
rect 1293 1053 1393 1069
rect 1293 1019 1309 1053
rect 1377 1019 1393 1053
rect 1293 972 1393 1019
rect 1451 1053 1551 1069
rect 1451 1019 1467 1053
rect 1535 1019 1551 1053
rect 1451 972 1551 1019
rect 1609 1053 1709 1069
rect 1609 1019 1625 1053
rect 1693 1019 1709 1053
rect 1609 972 1709 1019
rect 1767 1053 1867 1069
rect 1767 1019 1783 1053
rect 1851 1019 1867 1053
rect 1767 972 1867 1019
rect 1925 1053 2025 1069
rect 1925 1019 1941 1053
rect 2009 1019 2025 1053
rect 1925 972 2025 1019
rect 2083 1053 2183 1069
rect 2083 1019 2099 1053
rect 2167 1019 2183 1053
rect 2083 972 2183 1019
rect 2241 1053 2341 1069
rect 2241 1019 2257 1053
rect 2325 1019 2341 1053
rect 2241 972 2341 1019
rect 2399 1053 2499 1069
rect 2399 1019 2415 1053
rect 2483 1019 2499 1053
rect 2399 972 2499 1019
rect 2557 1053 2657 1069
rect 2557 1019 2573 1053
rect 2641 1019 2657 1053
rect 2557 972 2657 1019
rect 2715 1053 2815 1069
rect 2715 1019 2731 1053
rect 2799 1019 2815 1053
rect 2715 972 2815 1019
rect 2873 1053 2973 1069
rect 2873 1019 2889 1053
rect 2957 1019 2973 1053
rect 2873 972 2973 1019
rect 3031 1053 3131 1069
rect 3031 1019 3047 1053
rect 3115 1019 3131 1053
rect 3031 972 3131 1019
rect 3189 1053 3289 1069
rect 3189 1019 3205 1053
rect 3273 1019 3289 1053
rect 3189 972 3289 1019
rect 3347 1053 3447 1069
rect 3347 1019 3363 1053
rect 3431 1019 3447 1053
rect 3347 972 3447 1019
rect 3505 1053 3605 1069
rect 3505 1019 3521 1053
rect 3589 1019 3605 1053
rect 3505 972 3605 1019
rect 3663 1053 3763 1069
rect 3663 1019 3679 1053
rect 3747 1019 3763 1053
rect 3663 972 3763 1019
rect 3821 1053 3921 1069
rect 3821 1019 3837 1053
rect 3905 1019 3921 1053
rect 3821 972 3921 1019
rect 3979 1053 4079 1069
rect 3979 1019 3995 1053
rect 4063 1019 4079 1053
rect 3979 972 4079 1019
rect 4137 1053 4237 1069
rect 4137 1019 4153 1053
rect 4221 1019 4237 1053
rect 4137 972 4237 1019
rect 4295 1053 4395 1069
rect 4295 1019 4311 1053
rect 4379 1019 4395 1053
rect 4295 972 4395 1019
rect -4395 725 -4295 772
rect -4395 691 -4379 725
rect -4311 691 -4295 725
rect -4395 675 -4295 691
rect -4237 725 -4137 772
rect -4237 691 -4221 725
rect -4153 691 -4137 725
rect -4237 675 -4137 691
rect -4079 725 -3979 772
rect -4079 691 -4063 725
rect -3995 691 -3979 725
rect -4079 675 -3979 691
rect -3921 725 -3821 772
rect -3921 691 -3905 725
rect -3837 691 -3821 725
rect -3921 675 -3821 691
rect -3763 725 -3663 772
rect -3763 691 -3747 725
rect -3679 691 -3663 725
rect -3763 675 -3663 691
rect -3605 725 -3505 772
rect -3605 691 -3589 725
rect -3521 691 -3505 725
rect -3605 675 -3505 691
rect -3447 725 -3347 772
rect -3447 691 -3431 725
rect -3363 691 -3347 725
rect -3447 675 -3347 691
rect -3289 725 -3189 772
rect -3289 691 -3273 725
rect -3205 691 -3189 725
rect -3289 675 -3189 691
rect -3131 725 -3031 772
rect -3131 691 -3115 725
rect -3047 691 -3031 725
rect -3131 675 -3031 691
rect -2973 725 -2873 772
rect -2973 691 -2957 725
rect -2889 691 -2873 725
rect -2973 675 -2873 691
rect -2815 725 -2715 772
rect -2815 691 -2799 725
rect -2731 691 -2715 725
rect -2815 675 -2715 691
rect -2657 725 -2557 772
rect -2657 691 -2641 725
rect -2573 691 -2557 725
rect -2657 675 -2557 691
rect -2499 725 -2399 772
rect -2499 691 -2483 725
rect -2415 691 -2399 725
rect -2499 675 -2399 691
rect -2341 725 -2241 772
rect -2341 691 -2325 725
rect -2257 691 -2241 725
rect -2341 675 -2241 691
rect -2183 725 -2083 772
rect -2183 691 -2167 725
rect -2099 691 -2083 725
rect -2183 675 -2083 691
rect -2025 725 -1925 772
rect -2025 691 -2009 725
rect -1941 691 -1925 725
rect -2025 675 -1925 691
rect -1867 725 -1767 772
rect -1867 691 -1851 725
rect -1783 691 -1767 725
rect -1867 675 -1767 691
rect -1709 725 -1609 772
rect -1709 691 -1693 725
rect -1625 691 -1609 725
rect -1709 675 -1609 691
rect -1551 725 -1451 772
rect -1551 691 -1535 725
rect -1467 691 -1451 725
rect -1551 675 -1451 691
rect -1393 725 -1293 772
rect -1393 691 -1377 725
rect -1309 691 -1293 725
rect -1393 675 -1293 691
rect -1235 725 -1135 772
rect -1235 691 -1219 725
rect -1151 691 -1135 725
rect -1235 675 -1135 691
rect -1077 725 -977 772
rect -1077 691 -1061 725
rect -993 691 -977 725
rect -1077 675 -977 691
rect -919 725 -819 772
rect -919 691 -903 725
rect -835 691 -819 725
rect -919 675 -819 691
rect -761 725 -661 772
rect -761 691 -745 725
rect -677 691 -661 725
rect -761 675 -661 691
rect -603 725 -503 772
rect -603 691 -587 725
rect -519 691 -503 725
rect -603 675 -503 691
rect -445 725 -345 772
rect -445 691 -429 725
rect -361 691 -345 725
rect -445 675 -345 691
rect -287 725 -187 772
rect -287 691 -271 725
rect -203 691 -187 725
rect -287 675 -187 691
rect -129 725 -29 772
rect -129 691 -113 725
rect -45 691 -29 725
rect -129 675 -29 691
rect 29 725 129 772
rect 29 691 45 725
rect 113 691 129 725
rect 29 675 129 691
rect 187 725 287 772
rect 187 691 203 725
rect 271 691 287 725
rect 187 675 287 691
rect 345 725 445 772
rect 345 691 361 725
rect 429 691 445 725
rect 345 675 445 691
rect 503 725 603 772
rect 503 691 519 725
rect 587 691 603 725
rect 503 675 603 691
rect 661 725 761 772
rect 661 691 677 725
rect 745 691 761 725
rect 661 675 761 691
rect 819 725 919 772
rect 819 691 835 725
rect 903 691 919 725
rect 819 675 919 691
rect 977 725 1077 772
rect 977 691 993 725
rect 1061 691 1077 725
rect 977 675 1077 691
rect 1135 725 1235 772
rect 1135 691 1151 725
rect 1219 691 1235 725
rect 1135 675 1235 691
rect 1293 725 1393 772
rect 1293 691 1309 725
rect 1377 691 1393 725
rect 1293 675 1393 691
rect 1451 725 1551 772
rect 1451 691 1467 725
rect 1535 691 1551 725
rect 1451 675 1551 691
rect 1609 725 1709 772
rect 1609 691 1625 725
rect 1693 691 1709 725
rect 1609 675 1709 691
rect 1767 725 1867 772
rect 1767 691 1783 725
rect 1851 691 1867 725
rect 1767 675 1867 691
rect 1925 725 2025 772
rect 1925 691 1941 725
rect 2009 691 2025 725
rect 1925 675 2025 691
rect 2083 725 2183 772
rect 2083 691 2099 725
rect 2167 691 2183 725
rect 2083 675 2183 691
rect 2241 725 2341 772
rect 2241 691 2257 725
rect 2325 691 2341 725
rect 2241 675 2341 691
rect 2399 725 2499 772
rect 2399 691 2415 725
rect 2483 691 2499 725
rect 2399 675 2499 691
rect 2557 725 2657 772
rect 2557 691 2573 725
rect 2641 691 2657 725
rect 2557 675 2657 691
rect 2715 725 2815 772
rect 2715 691 2731 725
rect 2799 691 2815 725
rect 2715 675 2815 691
rect 2873 725 2973 772
rect 2873 691 2889 725
rect 2957 691 2973 725
rect 2873 675 2973 691
rect 3031 725 3131 772
rect 3031 691 3047 725
rect 3115 691 3131 725
rect 3031 675 3131 691
rect 3189 725 3289 772
rect 3189 691 3205 725
rect 3273 691 3289 725
rect 3189 675 3289 691
rect 3347 725 3447 772
rect 3347 691 3363 725
rect 3431 691 3447 725
rect 3347 675 3447 691
rect 3505 725 3605 772
rect 3505 691 3521 725
rect 3589 691 3605 725
rect 3505 675 3605 691
rect 3663 725 3763 772
rect 3663 691 3679 725
rect 3747 691 3763 725
rect 3663 675 3763 691
rect 3821 725 3921 772
rect 3821 691 3837 725
rect 3905 691 3921 725
rect 3821 675 3921 691
rect 3979 725 4079 772
rect 3979 691 3995 725
rect 4063 691 4079 725
rect 3979 675 4079 691
rect 4137 725 4237 772
rect 4137 691 4153 725
rect 4221 691 4237 725
rect 4137 675 4237 691
rect 4295 725 4395 772
rect 4295 691 4311 725
rect 4379 691 4395 725
rect 4295 675 4395 691
rect -4395 617 -4295 633
rect -4395 583 -4379 617
rect -4311 583 -4295 617
rect -4395 536 -4295 583
rect -4237 617 -4137 633
rect -4237 583 -4221 617
rect -4153 583 -4137 617
rect -4237 536 -4137 583
rect -4079 617 -3979 633
rect -4079 583 -4063 617
rect -3995 583 -3979 617
rect -4079 536 -3979 583
rect -3921 617 -3821 633
rect -3921 583 -3905 617
rect -3837 583 -3821 617
rect -3921 536 -3821 583
rect -3763 617 -3663 633
rect -3763 583 -3747 617
rect -3679 583 -3663 617
rect -3763 536 -3663 583
rect -3605 617 -3505 633
rect -3605 583 -3589 617
rect -3521 583 -3505 617
rect -3605 536 -3505 583
rect -3447 617 -3347 633
rect -3447 583 -3431 617
rect -3363 583 -3347 617
rect -3447 536 -3347 583
rect -3289 617 -3189 633
rect -3289 583 -3273 617
rect -3205 583 -3189 617
rect -3289 536 -3189 583
rect -3131 617 -3031 633
rect -3131 583 -3115 617
rect -3047 583 -3031 617
rect -3131 536 -3031 583
rect -2973 617 -2873 633
rect -2973 583 -2957 617
rect -2889 583 -2873 617
rect -2973 536 -2873 583
rect -2815 617 -2715 633
rect -2815 583 -2799 617
rect -2731 583 -2715 617
rect -2815 536 -2715 583
rect -2657 617 -2557 633
rect -2657 583 -2641 617
rect -2573 583 -2557 617
rect -2657 536 -2557 583
rect -2499 617 -2399 633
rect -2499 583 -2483 617
rect -2415 583 -2399 617
rect -2499 536 -2399 583
rect -2341 617 -2241 633
rect -2341 583 -2325 617
rect -2257 583 -2241 617
rect -2341 536 -2241 583
rect -2183 617 -2083 633
rect -2183 583 -2167 617
rect -2099 583 -2083 617
rect -2183 536 -2083 583
rect -2025 617 -1925 633
rect -2025 583 -2009 617
rect -1941 583 -1925 617
rect -2025 536 -1925 583
rect -1867 617 -1767 633
rect -1867 583 -1851 617
rect -1783 583 -1767 617
rect -1867 536 -1767 583
rect -1709 617 -1609 633
rect -1709 583 -1693 617
rect -1625 583 -1609 617
rect -1709 536 -1609 583
rect -1551 617 -1451 633
rect -1551 583 -1535 617
rect -1467 583 -1451 617
rect -1551 536 -1451 583
rect -1393 617 -1293 633
rect -1393 583 -1377 617
rect -1309 583 -1293 617
rect -1393 536 -1293 583
rect -1235 617 -1135 633
rect -1235 583 -1219 617
rect -1151 583 -1135 617
rect -1235 536 -1135 583
rect -1077 617 -977 633
rect -1077 583 -1061 617
rect -993 583 -977 617
rect -1077 536 -977 583
rect -919 617 -819 633
rect -919 583 -903 617
rect -835 583 -819 617
rect -919 536 -819 583
rect -761 617 -661 633
rect -761 583 -745 617
rect -677 583 -661 617
rect -761 536 -661 583
rect -603 617 -503 633
rect -603 583 -587 617
rect -519 583 -503 617
rect -603 536 -503 583
rect -445 617 -345 633
rect -445 583 -429 617
rect -361 583 -345 617
rect -445 536 -345 583
rect -287 617 -187 633
rect -287 583 -271 617
rect -203 583 -187 617
rect -287 536 -187 583
rect -129 617 -29 633
rect -129 583 -113 617
rect -45 583 -29 617
rect -129 536 -29 583
rect 29 617 129 633
rect 29 583 45 617
rect 113 583 129 617
rect 29 536 129 583
rect 187 617 287 633
rect 187 583 203 617
rect 271 583 287 617
rect 187 536 287 583
rect 345 617 445 633
rect 345 583 361 617
rect 429 583 445 617
rect 345 536 445 583
rect 503 617 603 633
rect 503 583 519 617
rect 587 583 603 617
rect 503 536 603 583
rect 661 617 761 633
rect 661 583 677 617
rect 745 583 761 617
rect 661 536 761 583
rect 819 617 919 633
rect 819 583 835 617
rect 903 583 919 617
rect 819 536 919 583
rect 977 617 1077 633
rect 977 583 993 617
rect 1061 583 1077 617
rect 977 536 1077 583
rect 1135 617 1235 633
rect 1135 583 1151 617
rect 1219 583 1235 617
rect 1135 536 1235 583
rect 1293 617 1393 633
rect 1293 583 1309 617
rect 1377 583 1393 617
rect 1293 536 1393 583
rect 1451 617 1551 633
rect 1451 583 1467 617
rect 1535 583 1551 617
rect 1451 536 1551 583
rect 1609 617 1709 633
rect 1609 583 1625 617
rect 1693 583 1709 617
rect 1609 536 1709 583
rect 1767 617 1867 633
rect 1767 583 1783 617
rect 1851 583 1867 617
rect 1767 536 1867 583
rect 1925 617 2025 633
rect 1925 583 1941 617
rect 2009 583 2025 617
rect 1925 536 2025 583
rect 2083 617 2183 633
rect 2083 583 2099 617
rect 2167 583 2183 617
rect 2083 536 2183 583
rect 2241 617 2341 633
rect 2241 583 2257 617
rect 2325 583 2341 617
rect 2241 536 2341 583
rect 2399 617 2499 633
rect 2399 583 2415 617
rect 2483 583 2499 617
rect 2399 536 2499 583
rect 2557 617 2657 633
rect 2557 583 2573 617
rect 2641 583 2657 617
rect 2557 536 2657 583
rect 2715 617 2815 633
rect 2715 583 2731 617
rect 2799 583 2815 617
rect 2715 536 2815 583
rect 2873 617 2973 633
rect 2873 583 2889 617
rect 2957 583 2973 617
rect 2873 536 2973 583
rect 3031 617 3131 633
rect 3031 583 3047 617
rect 3115 583 3131 617
rect 3031 536 3131 583
rect 3189 617 3289 633
rect 3189 583 3205 617
rect 3273 583 3289 617
rect 3189 536 3289 583
rect 3347 617 3447 633
rect 3347 583 3363 617
rect 3431 583 3447 617
rect 3347 536 3447 583
rect 3505 617 3605 633
rect 3505 583 3521 617
rect 3589 583 3605 617
rect 3505 536 3605 583
rect 3663 617 3763 633
rect 3663 583 3679 617
rect 3747 583 3763 617
rect 3663 536 3763 583
rect 3821 617 3921 633
rect 3821 583 3837 617
rect 3905 583 3921 617
rect 3821 536 3921 583
rect 3979 617 4079 633
rect 3979 583 3995 617
rect 4063 583 4079 617
rect 3979 536 4079 583
rect 4137 617 4237 633
rect 4137 583 4153 617
rect 4221 583 4237 617
rect 4137 536 4237 583
rect 4295 617 4395 633
rect 4295 583 4311 617
rect 4379 583 4395 617
rect 4295 536 4395 583
rect -4395 289 -4295 336
rect -4395 255 -4379 289
rect -4311 255 -4295 289
rect -4395 239 -4295 255
rect -4237 289 -4137 336
rect -4237 255 -4221 289
rect -4153 255 -4137 289
rect -4237 239 -4137 255
rect -4079 289 -3979 336
rect -4079 255 -4063 289
rect -3995 255 -3979 289
rect -4079 239 -3979 255
rect -3921 289 -3821 336
rect -3921 255 -3905 289
rect -3837 255 -3821 289
rect -3921 239 -3821 255
rect -3763 289 -3663 336
rect -3763 255 -3747 289
rect -3679 255 -3663 289
rect -3763 239 -3663 255
rect -3605 289 -3505 336
rect -3605 255 -3589 289
rect -3521 255 -3505 289
rect -3605 239 -3505 255
rect -3447 289 -3347 336
rect -3447 255 -3431 289
rect -3363 255 -3347 289
rect -3447 239 -3347 255
rect -3289 289 -3189 336
rect -3289 255 -3273 289
rect -3205 255 -3189 289
rect -3289 239 -3189 255
rect -3131 289 -3031 336
rect -3131 255 -3115 289
rect -3047 255 -3031 289
rect -3131 239 -3031 255
rect -2973 289 -2873 336
rect -2973 255 -2957 289
rect -2889 255 -2873 289
rect -2973 239 -2873 255
rect -2815 289 -2715 336
rect -2815 255 -2799 289
rect -2731 255 -2715 289
rect -2815 239 -2715 255
rect -2657 289 -2557 336
rect -2657 255 -2641 289
rect -2573 255 -2557 289
rect -2657 239 -2557 255
rect -2499 289 -2399 336
rect -2499 255 -2483 289
rect -2415 255 -2399 289
rect -2499 239 -2399 255
rect -2341 289 -2241 336
rect -2341 255 -2325 289
rect -2257 255 -2241 289
rect -2341 239 -2241 255
rect -2183 289 -2083 336
rect -2183 255 -2167 289
rect -2099 255 -2083 289
rect -2183 239 -2083 255
rect -2025 289 -1925 336
rect -2025 255 -2009 289
rect -1941 255 -1925 289
rect -2025 239 -1925 255
rect -1867 289 -1767 336
rect -1867 255 -1851 289
rect -1783 255 -1767 289
rect -1867 239 -1767 255
rect -1709 289 -1609 336
rect -1709 255 -1693 289
rect -1625 255 -1609 289
rect -1709 239 -1609 255
rect -1551 289 -1451 336
rect -1551 255 -1535 289
rect -1467 255 -1451 289
rect -1551 239 -1451 255
rect -1393 289 -1293 336
rect -1393 255 -1377 289
rect -1309 255 -1293 289
rect -1393 239 -1293 255
rect -1235 289 -1135 336
rect -1235 255 -1219 289
rect -1151 255 -1135 289
rect -1235 239 -1135 255
rect -1077 289 -977 336
rect -1077 255 -1061 289
rect -993 255 -977 289
rect -1077 239 -977 255
rect -919 289 -819 336
rect -919 255 -903 289
rect -835 255 -819 289
rect -919 239 -819 255
rect -761 289 -661 336
rect -761 255 -745 289
rect -677 255 -661 289
rect -761 239 -661 255
rect -603 289 -503 336
rect -603 255 -587 289
rect -519 255 -503 289
rect -603 239 -503 255
rect -445 289 -345 336
rect -445 255 -429 289
rect -361 255 -345 289
rect -445 239 -345 255
rect -287 289 -187 336
rect -287 255 -271 289
rect -203 255 -187 289
rect -287 239 -187 255
rect -129 289 -29 336
rect -129 255 -113 289
rect -45 255 -29 289
rect -129 239 -29 255
rect 29 289 129 336
rect 29 255 45 289
rect 113 255 129 289
rect 29 239 129 255
rect 187 289 287 336
rect 187 255 203 289
rect 271 255 287 289
rect 187 239 287 255
rect 345 289 445 336
rect 345 255 361 289
rect 429 255 445 289
rect 345 239 445 255
rect 503 289 603 336
rect 503 255 519 289
rect 587 255 603 289
rect 503 239 603 255
rect 661 289 761 336
rect 661 255 677 289
rect 745 255 761 289
rect 661 239 761 255
rect 819 289 919 336
rect 819 255 835 289
rect 903 255 919 289
rect 819 239 919 255
rect 977 289 1077 336
rect 977 255 993 289
rect 1061 255 1077 289
rect 977 239 1077 255
rect 1135 289 1235 336
rect 1135 255 1151 289
rect 1219 255 1235 289
rect 1135 239 1235 255
rect 1293 289 1393 336
rect 1293 255 1309 289
rect 1377 255 1393 289
rect 1293 239 1393 255
rect 1451 289 1551 336
rect 1451 255 1467 289
rect 1535 255 1551 289
rect 1451 239 1551 255
rect 1609 289 1709 336
rect 1609 255 1625 289
rect 1693 255 1709 289
rect 1609 239 1709 255
rect 1767 289 1867 336
rect 1767 255 1783 289
rect 1851 255 1867 289
rect 1767 239 1867 255
rect 1925 289 2025 336
rect 1925 255 1941 289
rect 2009 255 2025 289
rect 1925 239 2025 255
rect 2083 289 2183 336
rect 2083 255 2099 289
rect 2167 255 2183 289
rect 2083 239 2183 255
rect 2241 289 2341 336
rect 2241 255 2257 289
rect 2325 255 2341 289
rect 2241 239 2341 255
rect 2399 289 2499 336
rect 2399 255 2415 289
rect 2483 255 2499 289
rect 2399 239 2499 255
rect 2557 289 2657 336
rect 2557 255 2573 289
rect 2641 255 2657 289
rect 2557 239 2657 255
rect 2715 289 2815 336
rect 2715 255 2731 289
rect 2799 255 2815 289
rect 2715 239 2815 255
rect 2873 289 2973 336
rect 2873 255 2889 289
rect 2957 255 2973 289
rect 2873 239 2973 255
rect 3031 289 3131 336
rect 3031 255 3047 289
rect 3115 255 3131 289
rect 3031 239 3131 255
rect 3189 289 3289 336
rect 3189 255 3205 289
rect 3273 255 3289 289
rect 3189 239 3289 255
rect 3347 289 3447 336
rect 3347 255 3363 289
rect 3431 255 3447 289
rect 3347 239 3447 255
rect 3505 289 3605 336
rect 3505 255 3521 289
rect 3589 255 3605 289
rect 3505 239 3605 255
rect 3663 289 3763 336
rect 3663 255 3679 289
rect 3747 255 3763 289
rect 3663 239 3763 255
rect 3821 289 3921 336
rect 3821 255 3837 289
rect 3905 255 3921 289
rect 3821 239 3921 255
rect 3979 289 4079 336
rect 3979 255 3995 289
rect 4063 255 4079 289
rect 3979 239 4079 255
rect 4137 289 4237 336
rect 4137 255 4153 289
rect 4221 255 4237 289
rect 4137 239 4237 255
rect 4295 289 4395 336
rect 4295 255 4311 289
rect 4379 255 4395 289
rect 4295 239 4395 255
rect -4395 181 -4295 197
rect -4395 147 -4379 181
rect -4311 147 -4295 181
rect -4395 100 -4295 147
rect -4237 181 -4137 197
rect -4237 147 -4221 181
rect -4153 147 -4137 181
rect -4237 100 -4137 147
rect -4079 181 -3979 197
rect -4079 147 -4063 181
rect -3995 147 -3979 181
rect -4079 100 -3979 147
rect -3921 181 -3821 197
rect -3921 147 -3905 181
rect -3837 147 -3821 181
rect -3921 100 -3821 147
rect -3763 181 -3663 197
rect -3763 147 -3747 181
rect -3679 147 -3663 181
rect -3763 100 -3663 147
rect -3605 181 -3505 197
rect -3605 147 -3589 181
rect -3521 147 -3505 181
rect -3605 100 -3505 147
rect -3447 181 -3347 197
rect -3447 147 -3431 181
rect -3363 147 -3347 181
rect -3447 100 -3347 147
rect -3289 181 -3189 197
rect -3289 147 -3273 181
rect -3205 147 -3189 181
rect -3289 100 -3189 147
rect -3131 181 -3031 197
rect -3131 147 -3115 181
rect -3047 147 -3031 181
rect -3131 100 -3031 147
rect -2973 181 -2873 197
rect -2973 147 -2957 181
rect -2889 147 -2873 181
rect -2973 100 -2873 147
rect -2815 181 -2715 197
rect -2815 147 -2799 181
rect -2731 147 -2715 181
rect -2815 100 -2715 147
rect -2657 181 -2557 197
rect -2657 147 -2641 181
rect -2573 147 -2557 181
rect -2657 100 -2557 147
rect -2499 181 -2399 197
rect -2499 147 -2483 181
rect -2415 147 -2399 181
rect -2499 100 -2399 147
rect -2341 181 -2241 197
rect -2341 147 -2325 181
rect -2257 147 -2241 181
rect -2341 100 -2241 147
rect -2183 181 -2083 197
rect -2183 147 -2167 181
rect -2099 147 -2083 181
rect -2183 100 -2083 147
rect -2025 181 -1925 197
rect -2025 147 -2009 181
rect -1941 147 -1925 181
rect -2025 100 -1925 147
rect -1867 181 -1767 197
rect -1867 147 -1851 181
rect -1783 147 -1767 181
rect -1867 100 -1767 147
rect -1709 181 -1609 197
rect -1709 147 -1693 181
rect -1625 147 -1609 181
rect -1709 100 -1609 147
rect -1551 181 -1451 197
rect -1551 147 -1535 181
rect -1467 147 -1451 181
rect -1551 100 -1451 147
rect -1393 181 -1293 197
rect -1393 147 -1377 181
rect -1309 147 -1293 181
rect -1393 100 -1293 147
rect -1235 181 -1135 197
rect -1235 147 -1219 181
rect -1151 147 -1135 181
rect -1235 100 -1135 147
rect -1077 181 -977 197
rect -1077 147 -1061 181
rect -993 147 -977 181
rect -1077 100 -977 147
rect -919 181 -819 197
rect -919 147 -903 181
rect -835 147 -819 181
rect -919 100 -819 147
rect -761 181 -661 197
rect -761 147 -745 181
rect -677 147 -661 181
rect -761 100 -661 147
rect -603 181 -503 197
rect -603 147 -587 181
rect -519 147 -503 181
rect -603 100 -503 147
rect -445 181 -345 197
rect -445 147 -429 181
rect -361 147 -345 181
rect -445 100 -345 147
rect -287 181 -187 197
rect -287 147 -271 181
rect -203 147 -187 181
rect -287 100 -187 147
rect -129 181 -29 197
rect -129 147 -113 181
rect -45 147 -29 181
rect -129 100 -29 147
rect 29 181 129 197
rect 29 147 45 181
rect 113 147 129 181
rect 29 100 129 147
rect 187 181 287 197
rect 187 147 203 181
rect 271 147 287 181
rect 187 100 287 147
rect 345 181 445 197
rect 345 147 361 181
rect 429 147 445 181
rect 345 100 445 147
rect 503 181 603 197
rect 503 147 519 181
rect 587 147 603 181
rect 503 100 603 147
rect 661 181 761 197
rect 661 147 677 181
rect 745 147 761 181
rect 661 100 761 147
rect 819 181 919 197
rect 819 147 835 181
rect 903 147 919 181
rect 819 100 919 147
rect 977 181 1077 197
rect 977 147 993 181
rect 1061 147 1077 181
rect 977 100 1077 147
rect 1135 181 1235 197
rect 1135 147 1151 181
rect 1219 147 1235 181
rect 1135 100 1235 147
rect 1293 181 1393 197
rect 1293 147 1309 181
rect 1377 147 1393 181
rect 1293 100 1393 147
rect 1451 181 1551 197
rect 1451 147 1467 181
rect 1535 147 1551 181
rect 1451 100 1551 147
rect 1609 181 1709 197
rect 1609 147 1625 181
rect 1693 147 1709 181
rect 1609 100 1709 147
rect 1767 181 1867 197
rect 1767 147 1783 181
rect 1851 147 1867 181
rect 1767 100 1867 147
rect 1925 181 2025 197
rect 1925 147 1941 181
rect 2009 147 2025 181
rect 1925 100 2025 147
rect 2083 181 2183 197
rect 2083 147 2099 181
rect 2167 147 2183 181
rect 2083 100 2183 147
rect 2241 181 2341 197
rect 2241 147 2257 181
rect 2325 147 2341 181
rect 2241 100 2341 147
rect 2399 181 2499 197
rect 2399 147 2415 181
rect 2483 147 2499 181
rect 2399 100 2499 147
rect 2557 181 2657 197
rect 2557 147 2573 181
rect 2641 147 2657 181
rect 2557 100 2657 147
rect 2715 181 2815 197
rect 2715 147 2731 181
rect 2799 147 2815 181
rect 2715 100 2815 147
rect 2873 181 2973 197
rect 2873 147 2889 181
rect 2957 147 2973 181
rect 2873 100 2973 147
rect 3031 181 3131 197
rect 3031 147 3047 181
rect 3115 147 3131 181
rect 3031 100 3131 147
rect 3189 181 3289 197
rect 3189 147 3205 181
rect 3273 147 3289 181
rect 3189 100 3289 147
rect 3347 181 3447 197
rect 3347 147 3363 181
rect 3431 147 3447 181
rect 3347 100 3447 147
rect 3505 181 3605 197
rect 3505 147 3521 181
rect 3589 147 3605 181
rect 3505 100 3605 147
rect 3663 181 3763 197
rect 3663 147 3679 181
rect 3747 147 3763 181
rect 3663 100 3763 147
rect 3821 181 3921 197
rect 3821 147 3837 181
rect 3905 147 3921 181
rect 3821 100 3921 147
rect 3979 181 4079 197
rect 3979 147 3995 181
rect 4063 147 4079 181
rect 3979 100 4079 147
rect 4137 181 4237 197
rect 4137 147 4153 181
rect 4221 147 4237 181
rect 4137 100 4237 147
rect 4295 181 4395 197
rect 4295 147 4311 181
rect 4379 147 4395 181
rect 4295 100 4395 147
rect -4395 -147 -4295 -100
rect -4395 -181 -4379 -147
rect -4311 -181 -4295 -147
rect -4395 -197 -4295 -181
rect -4237 -147 -4137 -100
rect -4237 -181 -4221 -147
rect -4153 -181 -4137 -147
rect -4237 -197 -4137 -181
rect -4079 -147 -3979 -100
rect -4079 -181 -4063 -147
rect -3995 -181 -3979 -147
rect -4079 -197 -3979 -181
rect -3921 -147 -3821 -100
rect -3921 -181 -3905 -147
rect -3837 -181 -3821 -147
rect -3921 -197 -3821 -181
rect -3763 -147 -3663 -100
rect -3763 -181 -3747 -147
rect -3679 -181 -3663 -147
rect -3763 -197 -3663 -181
rect -3605 -147 -3505 -100
rect -3605 -181 -3589 -147
rect -3521 -181 -3505 -147
rect -3605 -197 -3505 -181
rect -3447 -147 -3347 -100
rect -3447 -181 -3431 -147
rect -3363 -181 -3347 -147
rect -3447 -197 -3347 -181
rect -3289 -147 -3189 -100
rect -3289 -181 -3273 -147
rect -3205 -181 -3189 -147
rect -3289 -197 -3189 -181
rect -3131 -147 -3031 -100
rect -3131 -181 -3115 -147
rect -3047 -181 -3031 -147
rect -3131 -197 -3031 -181
rect -2973 -147 -2873 -100
rect -2973 -181 -2957 -147
rect -2889 -181 -2873 -147
rect -2973 -197 -2873 -181
rect -2815 -147 -2715 -100
rect -2815 -181 -2799 -147
rect -2731 -181 -2715 -147
rect -2815 -197 -2715 -181
rect -2657 -147 -2557 -100
rect -2657 -181 -2641 -147
rect -2573 -181 -2557 -147
rect -2657 -197 -2557 -181
rect -2499 -147 -2399 -100
rect -2499 -181 -2483 -147
rect -2415 -181 -2399 -147
rect -2499 -197 -2399 -181
rect -2341 -147 -2241 -100
rect -2341 -181 -2325 -147
rect -2257 -181 -2241 -147
rect -2341 -197 -2241 -181
rect -2183 -147 -2083 -100
rect -2183 -181 -2167 -147
rect -2099 -181 -2083 -147
rect -2183 -197 -2083 -181
rect -2025 -147 -1925 -100
rect -2025 -181 -2009 -147
rect -1941 -181 -1925 -147
rect -2025 -197 -1925 -181
rect -1867 -147 -1767 -100
rect -1867 -181 -1851 -147
rect -1783 -181 -1767 -147
rect -1867 -197 -1767 -181
rect -1709 -147 -1609 -100
rect -1709 -181 -1693 -147
rect -1625 -181 -1609 -147
rect -1709 -197 -1609 -181
rect -1551 -147 -1451 -100
rect -1551 -181 -1535 -147
rect -1467 -181 -1451 -147
rect -1551 -197 -1451 -181
rect -1393 -147 -1293 -100
rect -1393 -181 -1377 -147
rect -1309 -181 -1293 -147
rect -1393 -197 -1293 -181
rect -1235 -147 -1135 -100
rect -1235 -181 -1219 -147
rect -1151 -181 -1135 -147
rect -1235 -197 -1135 -181
rect -1077 -147 -977 -100
rect -1077 -181 -1061 -147
rect -993 -181 -977 -147
rect -1077 -197 -977 -181
rect -919 -147 -819 -100
rect -919 -181 -903 -147
rect -835 -181 -819 -147
rect -919 -197 -819 -181
rect -761 -147 -661 -100
rect -761 -181 -745 -147
rect -677 -181 -661 -147
rect -761 -197 -661 -181
rect -603 -147 -503 -100
rect -603 -181 -587 -147
rect -519 -181 -503 -147
rect -603 -197 -503 -181
rect -445 -147 -345 -100
rect -445 -181 -429 -147
rect -361 -181 -345 -147
rect -445 -197 -345 -181
rect -287 -147 -187 -100
rect -287 -181 -271 -147
rect -203 -181 -187 -147
rect -287 -197 -187 -181
rect -129 -147 -29 -100
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect -129 -197 -29 -181
rect 29 -147 129 -100
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 29 -197 129 -181
rect 187 -147 287 -100
rect 187 -181 203 -147
rect 271 -181 287 -147
rect 187 -197 287 -181
rect 345 -147 445 -100
rect 345 -181 361 -147
rect 429 -181 445 -147
rect 345 -197 445 -181
rect 503 -147 603 -100
rect 503 -181 519 -147
rect 587 -181 603 -147
rect 503 -197 603 -181
rect 661 -147 761 -100
rect 661 -181 677 -147
rect 745 -181 761 -147
rect 661 -197 761 -181
rect 819 -147 919 -100
rect 819 -181 835 -147
rect 903 -181 919 -147
rect 819 -197 919 -181
rect 977 -147 1077 -100
rect 977 -181 993 -147
rect 1061 -181 1077 -147
rect 977 -197 1077 -181
rect 1135 -147 1235 -100
rect 1135 -181 1151 -147
rect 1219 -181 1235 -147
rect 1135 -197 1235 -181
rect 1293 -147 1393 -100
rect 1293 -181 1309 -147
rect 1377 -181 1393 -147
rect 1293 -197 1393 -181
rect 1451 -147 1551 -100
rect 1451 -181 1467 -147
rect 1535 -181 1551 -147
rect 1451 -197 1551 -181
rect 1609 -147 1709 -100
rect 1609 -181 1625 -147
rect 1693 -181 1709 -147
rect 1609 -197 1709 -181
rect 1767 -147 1867 -100
rect 1767 -181 1783 -147
rect 1851 -181 1867 -147
rect 1767 -197 1867 -181
rect 1925 -147 2025 -100
rect 1925 -181 1941 -147
rect 2009 -181 2025 -147
rect 1925 -197 2025 -181
rect 2083 -147 2183 -100
rect 2083 -181 2099 -147
rect 2167 -181 2183 -147
rect 2083 -197 2183 -181
rect 2241 -147 2341 -100
rect 2241 -181 2257 -147
rect 2325 -181 2341 -147
rect 2241 -197 2341 -181
rect 2399 -147 2499 -100
rect 2399 -181 2415 -147
rect 2483 -181 2499 -147
rect 2399 -197 2499 -181
rect 2557 -147 2657 -100
rect 2557 -181 2573 -147
rect 2641 -181 2657 -147
rect 2557 -197 2657 -181
rect 2715 -147 2815 -100
rect 2715 -181 2731 -147
rect 2799 -181 2815 -147
rect 2715 -197 2815 -181
rect 2873 -147 2973 -100
rect 2873 -181 2889 -147
rect 2957 -181 2973 -147
rect 2873 -197 2973 -181
rect 3031 -147 3131 -100
rect 3031 -181 3047 -147
rect 3115 -181 3131 -147
rect 3031 -197 3131 -181
rect 3189 -147 3289 -100
rect 3189 -181 3205 -147
rect 3273 -181 3289 -147
rect 3189 -197 3289 -181
rect 3347 -147 3447 -100
rect 3347 -181 3363 -147
rect 3431 -181 3447 -147
rect 3347 -197 3447 -181
rect 3505 -147 3605 -100
rect 3505 -181 3521 -147
rect 3589 -181 3605 -147
rect 3505 -197 3605 -181
rect 3663 -147 3763 -100
rect 3663 -181 3679 -147
rect 3747 -181 3763 -147
rect 3663 -197 3763 -181
rect 3821 -147 3921 -100
rect 3821 -181 3837 -147
rect 3905 -181 3921 -147
rect 3821 -197 3921 -181
rect 3979 -147 4079 -100
rect 3979 -181 3995 -147
rect 4063 -181 4079 -147
rect 3979 -197 4079 -181
rect 4137 -147 4237 -100
rect 4137 -181 4153 -147
rect 4221 -181 4237 -147
rect 4137 -197 4237 -181
rect 4295 -147 4395 -100
rect 4295 -181 4311 -147
rect 4379 -181 4395 -147
rect 4295 -197 4395 -181
rect -4395 -255 -4295 -239
rect -4395 -289 -4379 -255
rect -4311 -289 -4295 -255
rect -4395 -336 -4295 -289
rect -4237 -255 -4137 -239
rect -4237 -289 -4221 -255
rect -4153 -289 -4137 -255
rect -4237 -336 -4137 -289
rect -4079 -255 -3979 -239
rect -4079 -289 -4063 -255
rect -3995 -289 -3979 -255
rect -4079 -336 -3979 -289
rect -3921 -255 -3821 -239
rect -3921 -289 -3905 -255
rect -3837 -289 -3821 -255
rect -3921 -336 -3821 -289
rect -3763 -255 -3663 -239
rect -3763 -289 -3747 -255
rect -3679 -289 -3663 -255
rect -3763 -336 -3663 -289
rect -3605 -255 -3505 -239
rect -3605 -289 -3589 -255
rect -3521 -289 -3505 -255
rect -3605 -336 -3505 -289
rect -3447 -255 -3347 -239
rect -3447 -289 -3431 -255
rect -3363 -289 -3347 -255
rect -3447 -336 -3347 -289
rect -3289 -255 -3189 -239
rect -3289 -289 -3273 -255
rect -3205 -289 -3189 -255
rect -3289 -336 -3189 -289
rect -3131 -255 -3031 -239
rect -3131 -289 -3115 -255
rect -3047 -289 -3031 -255
rect -3131 -336 -3031 -289
rect -2973 -255 -2873 -239
rect -2973 -289 -2957 -255
rect -2889 -289 -2873 -255
rect -2973 -336 -2873 -289
rect -2815 -255 -2715 -239
rect -2815 -289 -2799 -255
rect -2731 -289 -2715 -255
rect -2815 -336 -2715 -289
rect -2657 -255 -2557 -239
rect -2657 -289 -2641 -255
rect -2573 -289 -2557 -255
rect -2657 -336 -2557 -289
rect -2499 -255 -2399 -239
rect -2499 -289 -2483 -255
rect -2415 -289 -2399 -255
rect -2499 -336 -2399 -289
rect -2341 -255 -2241 -239
rect -2341 -289 -2325 -255
rect -2257 -289 -2241 -255
rect -2341 -336 -2241 -289
rect -2183 -255 -2083 -239
rect -2183 -289 -2167 -255
rect -2099 -289 -2083 -255
rect -2183 -336 -2083 -289
rect -2025 -255 -1925 -239
rect -2025 -289 -2009 -255
rect -1941 -289 -1925 -255
rect -2025 -336 -1925 -289
rect -1867 -255 -1767 -239
rect -1867 -289 -1851 -255
rect -1783 -289 -1767 -255
rect -1867 -336 -1767 -289
rect -1709 -255 -1609 -239
rect -1709 -289 -1693 -255
rect -1625 -289 -1609 -255
rect -1709 -336 -1609 -289
rect -1551 -255 -1451 -239
rect -1551 -289 -1535 -255
rect -1467 -289 -1451 -255
rect -1551 -336 -1451 -289
rect -1393 -255 -1293 -239
rect -1393 -289 -1377 -255
rect -1309 -289 -1293 -255
rect -1393 -336 -1293 -289
rect -1235 -255 -1135 -239
rect -1235 -289 -1219 -255
rect -1151 -289 -1135 -255
rect -1235 -336 -1135 -289
rect -1077 -255 -977 -239
rect -1077 -289 -1061 -255
rect -993 -289 -977 -255
rect -1077 -336 -977 -289
rect -919 -255 -819 -239
rect -919 -289 -903 -255
rect -835 -289 -819 -255
rect -919 -336 -819 -289
rect -761 -255 -661 -239
rect -761 -289 -745 -255
rect -677 -289 -661 -255
rect -761 -336 -661 -289
rect -603 -255 -503 -239
rect -603 -289 -587 -255
rect -519 -289 -503 -255
rect -603 -336 -503 -289
rect -445 -255 -345 -239
rect -445 -289 -429 -255
rect -361 -289 -345 -255
rect -445 -336 -345 -289
rect -287 -255 -187 -239
rect -287 -289 -271 -255
rect -203 -289 -187 -255
rect -287 -336 -187 -289
rect -129 -255 -29 -239
rect -129 -289 -113 -255
rect -45 -289 -29 -255
rect -129 -336 -29 -289
rect 29 -255 129 -239
rect 29 -289 45 -255
rect 113 -289 129 -255
rect 29 -336 129 -289
rect 187 -255 287 -239
rect 187 -289 203 -255
rect 271 -289 287 -255
rect 187 -336 287 -289
rect 345 -255 445 -239
rect 345 -289 361 -255
rect 429 -289 445 -255
rect 345 -336 445 -289
rect 503 -255 603 -239
rect 503 -289 519 -255
rect 587 -289 603 -255
rect 503 -336 603 -289
rect 661 -255 761 -239
rect 661 -289 677 -255
rect 745 -289 761 -255
rect 661 -336 761 -289
rect 819 -255 919 -239
rect 819 -289 835 -255
rect 903 -289 919 -255
rect 819 -336 919 -289
rect 977 -255 1077 -239
rect 977 -289 993 -255
rect 1061 -289 1077 -255
rect 977 -336 1077 -289
rect 1135 -255 1235 -239
rect 1135 -289 1151 -255
rect 1219 -289 1235 -255
rect 1135 -336 1235 -289
rect 1293 -255 1393 -239
rect 1293 -289 1309 -255
rect 1377 -289 1393 -255
rect 1293 -336 1393 -289
rect 1451 -255 1551 -239
rect 1451 -289 1467 -255
rect 1535 -289 1551 -255
rect 1451 -336 1551 -289
rect 1609 -255 1709 -239
rect 1609 -289 1625 -255
rect 1693 -289 1709 -255
rect 1609 -336 1709 -289
rect 1767 -255 1867 -239
rect 1767 -289 1783 -255
rect 1851 -289 1867 -255
rect 1767 -336 1867 -289
rect 1925 -255 2025 -239
rect 1925 -289 1941 -255
rect 2009 -289 2025 -255
rect 1925 -336 2025 -289
rect 2083 -255 2183 -239
rect 2083 -289 2099 -255
rect 2167 -289 2183 -255
rect 2083 -336 2183 -289
rect 2241 -255 2341 -239
rect 2241 -289 2257 -255
rect 2325 -289 2341 -255
rect 2241 -336 2341 -289
rect 2399 -255 2499 -239
rect 2399 -289 2415 -255
rect 2483 -289 2499 -255
rect 2399 -336 2499 -289
rect 2557 -255 2657 -239
rect 2557 -289 2573 -255
rect 2641 -289 2657 -255
rect 2557 -336 2657 -289
rect 2715 -255 2815 -239
rect 2715 -289 2731 -255
rect 2799 -289 2815 -255
rect 2715 -336 2815 -289
rect 2873 -255 2973 -239
rect 2873 -289 2889 -255
rect 2957 -289 2973 -255
rect 2873 -336 2973 -289
rect 3031 -255 3131 -239
rect 3031 -289 3047 -255
rect 3115 -289 3131 -255
rect 3031 -336 3131 -289
rect 3189 -255 3289 -239
rect 3189 -289 3205 -255
rect 3273 -289 3289 -255
rect 3189 -336 3289 -289
rect 3347 -255 3447 -239
rect 3347 -289 3363 -255
rect 3431 -289 3447 -255
rect 3347 -336 3447 -289
rect 3505 -255 3605 -239
rect 3505 -289 3521 -255
rect 3589 -289 3605 -255
rect 3505 -336 3605 -289
rect 3663 -255 3763 -239
rect 3663 -289 3679 -255
rect 3747 -289 3763 -255
rect 3663 -336 3763 -289
rect 3821 -255 3921 -239
rect 3821 -289 3837 -255
rect 3905 -289 3921 -255
rect 3821 -336 3921 -289
rect 3979 -255 4079 -239
rect 3979 -289 3995 -255
rect 4063 -289 4079 -255
rect 3979 -336 4079 -289
rect 4137 -255 4237 -239
rect 4137 -289 4153 -255
rect 4221 -289 4237 -255
rect 4137 -336 4237 -289
rect 4295 -255 4395 -239
rect 4295 -289 4311 -255
rect 4379 -289 4395 -255
rect 4295 -336 4395 -289
rect -4395 -583 -4295 -536
rect -4395 -617 -4379 -583
rect -4311 -617 -4295 -583
rect -4395 -633 -4295 -617
rect -4237 -583 -4137 -536
rect -4237 -617 -4221 -583
rect -4153 -617 -4137 -583
rect -4237 -633 -4137 -617
rect -4079 -583 -3979 -536
rect -4079 -617 -4063 -583
rect -3995 -617 -3979 -583
rect -4079 -633 -3979 -617
rect -3921 -583 -3821 -536
rect -3921 -617 -3905 -583
rect -3837 -617 -3821 -583
rect -3921 -633 -3821 -617
rect -3763 -583 -3663 -536
rect -3763 -617 -3747 -583
rect -3679 -617 -3663 -583
rect -3763 -633 -3663 -617
rect -3605 -583 -3505 -536
rect -3605 -617 -3589 -583
rect -3521 -617 -3505 -583
rect -3605 -633 -3505 -617
rect -3447 -583 -3347 -536
rect -3447 -617 -3431 -583
rect -3363 -617 -3347 -583
rect -3447 -633 -3347 -617
rect -3289 -583 -3189 -536
rect -3289 -617 -3273 -583
rect -3205 -617 -3189 -583
rect -3289 -633 -3189 -617
rect -3131 -583 -3031 -536
rect -3131 -617 -3115 -583
rect -3047 -617 -3031 -583
rect -3131 -633 -3031 -617
rect -2973 -583 -2873 -536
rect -2973 -617 -2957 -583
rect -2889 -617 -2873 -583
rect -2973 -633 -2873 -617
rect -2815 -583 -2715 -536
rect -2815 -617 -2799 -583
rect -2731 -617 -2715 -583
rect -2815 -633 -2715 -617
rect -2657 -583 -2557 -536
rect -2657 -617 -2641 -583
rect -2573 -617 -2557 -583
rect -2657 -633 -2557 -617
rect -2499 -583 -2399 -536
rect -2499 -617 -2483 -583
rect -2415 -617 -2399 -583
rect -2499 -633 -2399 -617
rect -2341 -583 -2241 -536
rect -2341 -617 -2325 -583
rect -2257 -617 -2241 -583
rect -2341 -633 -2241 -617
rect -2183 -583 -2083 -536
rect -2183 -617 -2167 -583
rect -2099 -617 -2083 -583
rect -2183 -633 -2083 -617
rect -2025 -583 -1925 -536
rect -2025 -617 -2009 -583
rect -1941 -617 -1925 -583
rect -2025 -633 -1925 -617
rect -1867 -583 -1767 -536
rect -1867 -617 -1851 -583
rect -1783 -617 -1767 -583
rect -1867 -633 -1767 -617
rect -1709 -583 -1609 -536
rect -1709 -617 -1693 -583
rect -1625 -617 -1609 -583
rect -1709 -633 -1609 -617
rect -1551 -583 -1451 -536
rect -1551 -617 -1535 -583
rect -1467 -617 -1451 -583
rect -1551 -633 -1451 -617
rect -1393 -583 -1293 -536
rect -1393 -617 -1377 -583
rect -1309 -617 -1293 -583
rect -1393 -633 -1293 -617
rect -1235 -583 -1135 -536
rect -1235 -617 -1219 -583
rect -1151 -617 -1135 -583
rect -1235 -633 -1135 -617
rect -1077 -583 -977 -536
rect -1077 -617 -1061 -583
rect -993 -617 -977 -583
rect -1077 -633 -977 -617
rect -919 -583 -819 -536
rect -919 -617 -903 -583
rect -835 -617 -819 -583
rect -919 -633 -819 -617
rect -761 -583 -661 -536
rect -761 -617 -745 -583
rect -677 -617 -661 -583
rect -761 -633 -661 -617
rect -603 -583 -503 -536
rect -603 -617 -587 -583
rect -519 -617 -503 -583
rect -603 -633 -503 -617
rect -445 -583 -345 -536
rect -445 -617 -429 -583
rect -361 -617 -345 -583
rect -445 -633 -345 -617
rect -287 -583 -187 -536
rect -287 -617 -271 -583
rect -203 -617 -187 -583
rect -287 -633 -187 -617
rect -129 -583 -29 -536
rect -129 -617 -113 -583
rect -45 -617 -29 -583
rect -129 -633 -29 -617
rect 29 -583 129 -536
rect 29 -617 45 -583
rect 113 -617 129 -583
rect 29 -633 129 -617
rect 187 -583 287 -536
rect 187 -617 203 -583
rect 271 -617 287 -583
rect 187 -633 287 -617
rect 345 -583 445 -536
rect 345 -617 361 -583
rect 429 -617 445 -583
rect 345 -633 445 -617
rect 503 -583 603 -536
rect 503 -617 519 -583
rect 587 -617 603 -583
rect 503 -633 603 -617
rect 661 -583 761 -536
rect 661 -617 677 -583
rect 745 -617 761 -583
rect 661 -633 761 -617
rect 819 -583 919 -536
rect 819 -617 835 -583
rect 903 -617 919 -583
rect 819 -633 919 -617
rect 977 -583 1077 -536
rect 977 -617 993 -583
rect 1061 -617 1077 -583
rect 977 -633 1077 -617
rect 1135 -583 1235 -536
rect 1135 -617 1151 -583
rect 1219 -617 1235 -583
rect 1135 -633 1235 -617
rect 1293 -583 1393 -536
rect 1293 -617 1309 -583
rect 1377 -617 1393 -583
rect 1293 -633 1393 -617
rect 1451 -583 1551 -536
rect 1451 -617 1467 -583
rect 1535 -617 1551 -583
rect 1451 -633 1551 -617
rect 1609 -583 1709 -536
rect 1609 -617 1625 -583
rect 1693 -617 1709 -583
rect 1609 -633 1709 -617
rect 1767 -583 1867 -536
rect 1767 -617 1783 -583
rect 1851 -617 1867 -583
rect 1767 -633 1867 -617
rect 1925 -583 2025 -536
rect 1925 -617 1941 -583
rect 2009 -617 2025 -583
rect 1925 -633 2025 -617
rect 2083 -583 2183 -536
rect 2083 -617 2099 -583
rect 2167 -617 2183 -583
rect 2083 -633 2183 -617
rect 2241 -583 2341 -536
rect 2241 -617 2257 -583
rect 2325 -617 2341 -583
rect 2241 -633 2341 -617
rect 2399 -583 2499 -536
rect 2399 -617 2415 -583
rect 2483 -617 2499 -583
rect 2399 -633 2499 -617
rect 2557 -583 2657 -536
rect 2557 -617 2573 -583
rect 2641 -617 2657 -583
rect 2557 -633 2657 -617
rect 2715 -583 2815 -536
rect 2715 -617 2731 -583
rect 2799 -617 2815 -583
rect 2715 -633 2815 -617
rect 2873 -583 2973 -536
rect 2873 -617 2889 -583
rect 2957 -617 2973 -583
rect 2873 -633 2973 -617
rect 3031 -583 3131 -536
rect 3031 -617 3047 -583
rect 3115 -617 3131 -583
rect 3031 -633 3131 -617
rect 3189 -583 3289 -536
rect 3189 -617 3205 -583
rect 3273 -617 3289 -583
rect 3189 -633 3289 -617
rect 3347 -583 3447 -536
rect 3347 -617 3363 -583
rect 3431 -617 3447 -583
rect 3347 -633 3447 -617
rect 3505 -583 3605 -536
rect 3505 -617 3521 -583
rect 3589 -617 3605 -583
rect 3505 -633 3605 -617
rect 3663 -583 3763 -536
rect 3663 -617 3679 -583
rect 3747 -617 3763 -583
rect 3663 -633 3763 -617
rect 3821 -583 3921 -536
rect 3821 -617 3837 -583
rect 3905 -617 3921 -583
rect 3821 -633 3921 -617
rect 3979 -583 4079 -536
rect 3979 -617 3995 -583
rect 4063 -617 4079 -583
rect 3979 -633 4079 -617
rect 4137 -583 4237 -536
rect 4137 -617 4153 -583
rect 4221 -617 4237 -583
rect 4137 -633 4237 -617
rect 4295 -583 4395 -536
rect 4295 -617 4311 -583
rect 4379 -617 4395 -583
rect 4295 -633 4395 -617
rect -4395 -691 -4295 -675
rect -4395 -725 -4379 -691
rect -4311 -725 -4295 -691
rect -4395 -772 -4295 -725
rect -4237 -691 -4137 -675
rect -4237 -725 -4221 -691
rect -4153 -725 -4137 -691
rect -4237 -772 -4137 -725
rect -4079 -691 -3979 -675
rect -4079 -725 -4063 -691
rect -3995 -725 -3979 -691
rect -4079 -772 -3979 -725
rect -3921 -691 -3821 -675
rect -3921 -725 -3905 -691
rect -3837 -725 -3821 -691
rect -3921 -772 -3821 -725
rect -3763 -691 -3663 -675
rect -3763 -725 -3747 -691
rect -3679 -725 -3663 -691
rect -3763 -772 -3663 -725
rect -3605 -691 -3505 -675
rect -3605 -725 -3589 -691
rect -3521 -725 -3505 -691
rect -3605 -772 -3505 -725
rect -3447 -691 -3347 -675
rect -3447 -725 -3431 -691
rect -3363 -725 -3347 -691
rect -3447 -772 -3347 -725
rect -3289 -691 -3189 -675
rect -3289 -725 -3273 -691
rect -3205 -725 -3189 -691
rect -3289 -772 -3189 -725
rect -3131 -691 -3031 -675
rect -3131 -725 -3115 -691
rect -3047 -725 -3031 -691
rect -3131 -772 -3031 -725
rect -2973 -691 -2873 -675
rect -2973 -725 -2957 -691
rect -2889 -725 -2873 -691
rect -2973 -772 -2873 -725
rect -2815 -691 -2715 -675
rect -2815 -725 -2799 -691
rect -2731 -725 -2715 -691
rect -2815 -772 -2715 -725
rect -2657 -691 -2557 -675
rect -2657 -725 -2641 -691
rect -2573 -725 -2557 -691
rect -2657 -772 -2557 -725
rect -2499 -691 -2399 -675
rect -2499 -725 -2483 -691
rect -2415 -725 -2399 -691
rect -2499 -772 -2399 -725
rect -2341 -691 -2241 -675
rect -2341 -725 -2325 -691
rect -2257 -725 -2241 -691
rect -2341 -772 -2241 -725
rect -2183 -691 -2083 -675
rect -2183 -725 -2167 -691
rect -2099 -725 -2083 -691
rect -2183 -772 -2083 -725
rect -2025 -691 -1925 -675
rect -2025 -725 -2009 -691
rect -1941 -725 -1925 -691
rect -2025 -772 -1925 -725
rect -1867 -691 -1767 -675
rect -1867 -725 -1851 -691
rect -1783 -725 -1767 -691
rect -1867 -772 -1767 -725
rect -1709 -691 -1609 -675
rect -1709 -725 -1693 -691
rect -1625 -725 -1609 -691
rect -1709 -772 -1609 -725
rect -1551 -691 -1451 -675
rect -1551 -725 -1535 -691
rect -1467 -725 -1451 -691
rect -1551 -772 -1451 -725
rect -1393 -691 -1293 -675
rect -1393 -725 -1377 -691
rect -1309 -725 -1293 -691
rect -1393 -772 -1293 -725
rect -1235 -691 -1135 -675
rect -1235 -725 -1219 -691
rect -1151 -725 -1135 -691
rect -1235 -772 -1135 -725
rect -1077 -691 -977 -675
rect -1077 -725 -1061 -691
rect -993 -725 -977 -691
rect -1077 -772 -977 -725
rect -919 -691 -819 -675
rect -919 -725 -903 -691
rect -835 -725 -819 -691
rect -919 -772 -819 -725
rect -761 -691 -661 -675
rect -761 -725 -745 -691
rect -677 -725 -661 -691
rect -761 -772 -661 -725
rect -603 -691 -503 -675
rect -603 -725 -587 -691
rect -519 -725 -503 -691
rect -603 -772 -503 -725
rect -445 -691 -345 -675
rect -445 -725 -429 -691
rect -361 -725 -345 -691
rect -445 -772 -345 -725
rect -287 -691 -187 -675
rect -287 -725 -271 -691
rect -203 -725 -187 -691
rect -287 -772 -187 -725
rect -129 -691 -29 -675
rect -129 -725 -113 -691
rect -45 -725 -29 -691
rect -129 -772 -29 -725
rect 29 -691 129 -675
rect 29 -725 45 -691
rect 113 -725 129 -691
rect 29 -772 129 -725
rect 187 -691 287 -675
rect 187 -725 203 -691
rect 271 -725 287 -691
rect 187 -772 287 -725
rect 345 -691 445 -675
rect 345 -725 361 -691
rect 429 -725 445 -691
rect 345 -772 445 -725
rect 503 -691 603 -675
rect 503 -725 519 -691
rect 587 -725 603 -691
rect 503 -772 603 -725
rect 661 -691 761 -675
rect 661 -725 677 -691
rect 745 -725 761 -691
rect 661 -772 761 -725
rect 819 -691 919 -675
rect 819 -725 835 -691
rect 903 -725 919 -691
rect 819 -772 919 -725
rect 977 -691 1077 -675
rect 977 -725 993 -691
rect 1061 -725 1077 -691
rect 977 -772 1077 -725
rect 1135 -691 1235 -675
rect 1135 -725 1151 -691
rect 1219 -725 1235 -691
rect 1135 -772 1235 -725
rect 1293 -691 1393 -675
rect 1293 -725 1309 -691
rect 1377 -725 1393 -691
rect 1293 -772 1393 -725
rect 1451 -691 1551 -675
rect 1451 -725 1467 -691
rect 1535 -725 1551 -691
rect 1451 -772 1551 -725
rect 1609 -691 1709 -675
rect 1609 -725 1625 -691
rect 1693 -725 1709 -691
rect 1609 -772 1709 -725
rect 1767 -691 1867 -675
rect 1767 -725 1783 -691
rect 1851 -725 1867 -691
rect 1767 -772 1867 -725
rect 1925 -691 2025 -675
rect 1925 -725 1941 -691
rect 2009 -725 2025 -691
rect 1925 -772 2025 -725
rect 2083 -691 2183 -675
rect 2083 -725 2099 -691
rect 2167 -725 2183 -691
rect 2083 -772 2183 -725
rect 2241 -691 2341 -675
rect 2241 -725 2257 -691
rect 2325 -725 2341 -691
rect 2241 -772 2341 -725
rect 2399 -691 2499 -675
rect 2399 -725 2415 -691
rect 2483 -725 2499 -691
rect 2399 -772 2499 -725
rect 2557 -691 2657 -675
rect 2557 -725 2573 -691
rect 2641 -725 2657 -691
rect 2557 -772 2657 -725
rect 2715 -691 2815 -675
rect 2715 -725 2731 -691
rect 2799 -725 2815 -691
rect 2715 -772 2815 -725
rect 2873 -691 2973 -675
rect 2873 -725 2889 -691
rect 2957 -725 2973 -691
rect 2873 -772 2973 -725
rect 3031 -691 3131 -675
rect 3031 -725 3047 -691
rect 3115 -725 3131 -691
rect 3031 -772 3131 -725
rect 3189 -691 3289 -675
rect 3189 -725 3205 -691
rect 3273 -725 3289 -691
rect 3189 -772 3289 -725
rect 3347 -691 3447 -675
rect 3347 -725 3363 -691
rect 3431 -725 3447 -691
rect 3347 -772 3447 -725
rect 3505 -691 3605 -675
rect 3505 -725 3521 -691
rect 3589 -725 3605 -691
rect 3505 -772 3605 -725
rect 3663 -691 3763 -675
rect 3663 -725 3679 -691
rect 3747 -725 3763 -691
rect 3663 -772 3763 -725
rect 3821 -691 3921 -675
rect 3821 -725 3837 -691
rect 3905 -725 3921 -691
rect 3821 -772 3921 -725
rect 3979 -691 4079 -675
rect 3979 -725 3995 -691
rect 4063 -725 4079 -691
rect 3979 -772 4079 -725
rect 4137 -691 4237 -675
rect 4137 -725 4153 -691
rect 4221 -725 4237 -691
rect 4137 -772 4237 -725
rect 4295 -691 4395 -675
rect 4295 -725 4311 -691
rect 4379 -725 4395 -691
rect 4295 -772 4395 -725
rect -4395 -1019 -4295 -972
rect -4395 -1053 -4379 -1019
rect -4311 -1053 -4295 -1019
rect -4395 -1069 -4295 -1053
rect -4237 -1019 -4137 -972
rect -4237 -1053 -4221 -1019
rect -4153 -1053 -4137 -1019
rect -4237 -1069 -4137 -1053
rect -4079 -1019 -3979 -972
rect -4079 -1053 -4063 -1019
rect -3995 -1053 -3979 -1019
rect -4079 -1069 -3979 -1053
rect -3921 -1019 -3821 -972
rect -3921 -1053 -3905 -1019
rect -3837 -1053 -3821 -1019
rect -3921 -1069 -3821 -1053
rect -3763 -1019 -3663 -972
rect -3763 -1053 -3747 -1019
rect -3679 -1053 -3663 -1019
rect -3763 -1069 -3663 -1053
rect -3605 -1019 -3505 -972
rect -3605 -1053 -3589 -1019
rect -3521 -1053 -3505 -1019
rect -3605 -1069 -3505 -1053
rect -3447 -1019 -3347 -972
rect -3447 -1053 -3431 -1019
rect -3363 -1053 -3347 -1019
rect -3447 -1069 -3347 -1053
rect -3289 -1019 -3189 -972
rect -3289 -1053 -3273 -1019
rect -3205 -1053 -3189 -1019
rect -3289 -1069 -3189 -1053
rect -3131 -1019 -3031 -972
rect -3131 -1053 -3115 -1019
rect -3047 -1053 -3031 -1019
rect -3131 -1069 -3031 -1053
rect -2973 -1019 -2873 -972
rect -2973 -1053 -2957 -1019
rect -2889 -1053 -2873 -1019
rect -2973 -1069 -2873 -1053
rect -2815 -1019 -2715 -972
rect -2815 -1053 -2799 -1019
rect -2731 -1053 -2715 -1019
rect -2815 -1069 -2715 -1053
rect -2657 -1019 -2557 -972
rect -2657 -1053 -2641 -1019
rect -2573 -1053 -2557 -1019
rect -2657 -1069 -2557 -1053
rect -2499 -1019 -2399 -972
rect -2499 -1053 -2483 -1019
rect -2415 -1053 -2399 -1019
rect -2499 -1069 -2399 -1053
rect -2341 -1019 -2241 -972
rect -2341 -1053 -2325 -1019
rect -2257 -1053 -2241 -1019
rect -2341 -1069 -2241 -1053
rect -2183 -1019 -2083 -972
rect -2183 -1053 -2167 -1019
rect -2099 -1053 -2083 -1019
rect -2183 -1069 -2083 -1053
rect -2025 -1019 -1925 -972
rect -2025 -1053 -2009 -1019
rect -1941 -1053 -1925 -1019
rect -2025 -1069 -1925 -1053
rect -1867 -1019 -1767 -972
rect -1867 -1053 -1851 -1019
rect -1783 -1053 -1767 -1019
rect -1867 -1069 -1767 -1053
rect -1709 -1019 -1609 -972
rect -1709 -1053 -1693 -1019
rect -1625 -1053 -1609 -1019
rect -1709 -1069 -1609 -1053
rect -1551 -1019 -1451 -972
rect -1551 -1053 -1535 -1019
rect -1467 -1053 -1451 -1019
rect -1551 -1069 -1451 -1053
rect -1393 -1019 -1293 -972
rect -1393 -1053 -1377 -1019
rect -1309 -1053 -1293 -1019
rect -1393 -1069 -1293 -1053
rect -1235 -1019 -1135 -972
rect -1235 -1053 -1219 -1019
rect -1151 -1053 -1135 -1019
rect -1235 -1069 -1135 -1053
rect -1077 -1019 -977 -972
rect -1077 -1053 -1061 -1019
rect -993 -1053 -977 -1019
rect -1077 -1069 -977 -1053
rect -919 -1019 -819 -972
rect -919 -1053 -903 -1019
rect -835 -1053 -819 -1019
rect -919 -1069 -819 -1053
rect -761 -1019 -661 -972
rect -761 -1053 -745 -1019
rect -677 -1053 -661 -1019
rect -761 -1069 -661 -1053
rect -603 -1019 -503 -972
rect -603 -1053 -587 -1019
rect -519 -1053 -503 -1019
rect -603 -1069 -503 -1053
rect -445 -1019 -345 -972
rect -445 -1053 -429 -1019
rect -361 -1053 -345 -1019
rect -445 -1069 -345 -1053
rect -287 -1019 -187 -972
rect -287 -1053 -271 -1019
rect -203 -1053 -187 -1019
rect -287 -1069 -187 -1053
rect -129 -1019 -29 -972
rect -129 -1053 -113 -1019
rect -45 -1053 -29 -1019
rect -129 -1069 -29 -1053
rect 29 -1019 129 -972
rect 29 -1053 45 -1019
rect 113 -1053 129 -1019
rect 29 -1069 129 -1053
rect 187 -1019 287 -972
rect 187 -1053 203 -1019
rect 271 -1053 287 -1019
rect 187 -1069 287 -1053
rect 345 -1019 445 -972
rect 345 -1053 361 -1019
rect 429 -1053 445 -1019
rect 345 -1069 445 -1053
rect 503 -1019 603 -972
rect 503 -1053 519 -1019
rect 587 -1053 603 -1019
rect 503 -1069 603 -1053
rect 661 -1019 761 -972
rect 661 -1053 677 -1019
rect 745 -1053 761 -1019
rect 661 -1069 761 -1053
rect 819 -1019 919 -972
rect 819 -1053 835 -1019
rect 903 -1053 919 -1019
rect 819 -1069 919 -1053
rect 977 -1019 1077 -972
rect 977 -1053 993 -1019
rect 1061 -1053 1077 -1019
rect 977 -1069 1077 -1053
rect 1135 -1019 1235 -972
rect 1135 -1053 1151 -1019
rect 1219 -1053 1235 -1019
rect 1135 -1069 1235 -1053
rect 1293 -1019 1393 -972
rect 1293 -1053 1309 -1019
rect 1377 -1053 1393 -1019
rect 1293 -1069 1393 -1053
rect 1451 -1019 1551 -972
rect 1451 -1053 1467 -1019
rect 1535 -1053 1551 -1019
rect 1451 -1069 1551 -1053
rect 1609 -1019 1709 -972
rect 1609 -1053 1625 -1019
rect 1693 -1053 1709 -1019
rect 1609 -1069 1709 -1053
rect 1767 -1019 1867 -972
rect 1767 -1053 1783 -1019
rect 1851 -1053 1867 -1019
rect 1767 -1069 1867 -1053
rect 1925 -1019 2025 -972
rect 1925 -1053 1941 -1019
rect 2009 -1053 2025 -1019
rect 1925 -1069 2025 -1053
rect 2083 -1019 2183 -972
rect 2083 -1053 2099 -1019
rect 2167 -1053 2183 -1019
rect 2083 -1069 2183 -1053
rect 2241 -1019 2341 -972
rect 2241 -1053 2257 -1019
rect 2325 -1053 2341 -1019
rect 2241 -1069 2341 -1053
rect 2399 -1019 2499 -972
rect 2399 -1053 2415 -1019
rect 2483 -1053 2499 -1019
rect 2399 -1069 2499 -1053
rect 2557 -1019 2657 -972
rect 2557 -1053 2573 -1019
rect 2641 -1053 2657 -1019
rect 2557 -1069 2657 -1053
rect 2715 -1019 2815 -972
rect 2715 -1053 2731 -1019
rect 2799 -1053 2815 -1019
rect 2715 -1069 2815 -1053
rect 2873 -1019 2973 -972
rect 2873 -1053 2889 -1019
rect 2957 -1053 2973 -1019
rect 2873 -1069 2973 -1053
rect 3031 -1019 3131 -972
rect 3031 -1053 3047 -1019
rect 3115 -1053 3131 -1019
rect 3031 -1069 3131 -1053
rect 3189 -1019 3289 -972
rect 3189 -1053 3205 -1019
rect 3273 -1053 3289 -1019
rect 3189 -1069 3289 -1053
rect 3347 -1019 3447 -972
rect 3347 -1053 3363 -1019
rect 3431 -1053 3447 -1019
rect 3347 -1069 3447 -1053
rect 3505 -1019 3605 -972
rect 3505 -1053 3521 -1019
rect 3589 -1053 3605 -1019
rect 3505 -1069 3605 -1053
rect 3663 -1019 3763 -972
rect 3663 -1053 3679 -1019
rect 3747 -1053 3763 -1019
rect 3663 -1069 3763 -1053
rect 3821 -1019 3921 -972
rect 3821 -1053 3837 -1019
rect 3905 -1053 3921 -1019
rect 3821 -1069 3921 -1053
rect 3979 -1019 4079 -972
rect 3979 -1053 3995 -1019
rect 4063 -1053 4079 -1019
rect 3979 -1069 4079 -1053
rect 4137 -1019 4237 -972
rect 4137 -1053 4153 -1019
rect 4221 -1053 4237 -1019
rect 4137 -1069 4237 -1053
rect 4295 -1019 4395 -972
rect 4295 -1053 4311 -1019
rect 4379 -1053 4395 -1019
rect 4295 -1069 4395 -1053
<< polycont >>
rect -4379 1019 -4311 1053
rect -4221 1019 -4153 1053
rect -4063 1019 -3995 1053
rect -3905 1019 -3837 1053
rect -3747 1019 -3679 1053
rect -3589 1019 -3521 1053
rect -3431 1019 -3363 1053
rect -3273 1019 -3205 1053
rect -3115 1019 -3047 1053
rect -2957 1019 -2889 1053
rect -2799 1019 -2731 1053
rect -2641 1019 -2573 1053
rect -2483 1019 -2415 1053
rect -2325 1019 -2257 1053
rect -2167 1019 -2099 1053
rect -2009 1019 -1941 1053
rect -1851 1019 -1783 1053
rect -1693 1019 -1625 1053
rect -1535 1019 -1467 1053
rect -1377 1019 -1309 1053
rect -1219 1019 -1151 1053
rect -1061 1019 -993 1053
rect -903 1019 -835 1053
rect -745 1019 -677 1053
rect -587 1019 -519 1053
rect -429 1019 -361 1053
rect -271 1019 -203 1053
rect -113 1019 -45 1053
rect 45 1019 113 1053
rect 203 1019 271 1053
rect 361 1019 429 1053
rect 519 1019 587 1053
rect 677 1019 745 1053
rect 835 1019 903 1053
rect 993 1019 1061 1053
rect 1151 1019 1219 1053
rect 1309 1019 1377 1053
rect 1467 1019 1535 1053
rect 1625 1019 1693 1053
rect 1783 1019 1851 1053
rect 1941 1019 2009 1053
rect 2099 1019 2167 1053
rect 2257 1019 2325 1053
rect 2415 1019 2483 1053
rect 2573 1019 2641 1053
rect 2731 1019 2799 1053
rect 2889 1019 2957 1053
rect 3047 1019 3115 1053
rect 3205 1019 3273 1053
rect 3363 1019 3431 1053
rect 3521 1019 3589 1053
rect 3679 1019 3747 1053
rect 3837 1019 3905 1053
rect 3995 1019 4063 1053
rect 4153 1019 4221 1053
rect 4311 1019 4379 1053
rect -4379 691 -4311 725
rect -4221 691 -4153 725
rect -4063 691 -3995 725
rect -3905 691 -3837 725
rect -3747 691 -3679 725
rect -3589 691 -3521 725
rect -3431 691 -3363 725
rect -3273 691 -3205 725
rect -3115 691 -3047 725
rect -2957 691 -2889 725
rect -2799 691 -2731 725
rect -2641 691 -2573 725
rect -2483 691 -2415 725
rect -2325 691 -2257 725
rect -2167 691 -2099 725
rect -2009 691 -1941 725
rect -1851 691 -1783 725
rect -1693 691 -1625 725
rect -1535 691 -1467 725
rect -1377 691 -1309 725
rect -1219 691 -1151 725
rect -1061 691 -993 725
rect -903 691 -835 725
rect -745 691 -677 725
rect -587 691 -519 725
rect -429 691 -361 725
rect -271 691 -203 725
rect -113 691 -45 725
rect 45 691 113 725
rect 203 691 271 725
rect 361 691 429 725
rect 519 691 587 725
rect 677 691 745 725
rect 835 691 903 725
rect 993 691 1061 725
rect 1151 691 1219 725
rect 1309 691 1377 725
rect 1467 691 1535 725
rect 1625 691 1693 725
rect 1783 691 1851 725
rect 1941 691 2009 725
rect 2099 691 2167 725
rect 2257 691 2325 725
rect 2415 691 2483 725
rect 2573 691 2641 725
rect 2731 691 2799 725
rect 2889 691 2957 725
rect 3047 691 3115 725
rect 3205 691 3273 725
rect 3363 691 3431 725
rect 3521 691 3589 725
rect 3679 691 3747 725
rect 3837 691 3905 725
rect 3995 691 4063 725
rect 4153 691 4221 725
rect 4311 691 4379 725
rect -4379 583 -4311 617
rect -4221 583 -4153 617
rect -4063 583 -3995 617
rect -3905 583 -3837 617
rect -3747 583 -3679 617
rect -3589 583 -3521 617
rect -3431 583 -3363 617
rect -3273 583 -3205 617
rect -3115 583 -3047 617
rect -2957 583 -2889 617
rect -2799 583 -2731 617
rect -2641 583 -2573 617
rect -2483 583 -2415 617
rect -2325 583 -2257 617
rect -2167 583 -2099 617
rect -2009 583 -1941 617
rect -1851 583 -1783 617
rect -1693 583 -1625 617
rect -1535 583 -1467 617
rect -1377 583 -1309 617
rect -1219 583 -1151 617
rect -1061 583 -993 617
rect -903 583 -835 617
rect -745 583 -677 617
rect -587 583 -519 617
rect -429 583 -361 617
rect -271 583 -203 617
rect -113 583 -45 617
rect 45 583 113 617
rect 203 583 271 617
rect 361 583 429 617
rect 519 583 587 617
rect 677 583 745 617
rect 835 583 903 617
rect 993 583 1061 617
rect 1151 583 1219 617
rect 1309 583 1377 617
rect 1467 583 1535 617
rect 1625 583 1693 617
rect 1783 583 1851 617
rect 1941 583 2009 617
rect 2099 583 2167 617
rect 2257 583 2325 617
rect 2415 583 2483 617
rect 2573 583 2641 617
rect 2731 583 2799 617
rect 2889 583 2957 617
rect 3047 583 3115 617
rect 3205 583 3273 617
rect 3363 583 3431 617
rect 3521 583 3589 617
rect 3679 583 3747 617
rect 3837 583 3905 617
rect 3995 583 4063 617
rect 4153 583 4221 617
rect 4311 583 4379 617
rect -4379 255 -4311 289
rect -4221 255 -4153 289
rect -4063 255 -3995 289
rect -3905 255 -3837 289
rect -3747 255 -3679 289
rect -3589 255 -3521 289
rect -3431 255 -3363 289
rect -3273 255 -3205 289
rect -3115 255 -3047 289
rect -2957 255 -2889 289
rect -2799 255 -2731 289
rect -2641 255 -2573 289
rect -2483 255 -2415 289
rect -2325 255 -2257 289
rect -2167 255 -2099 289
rect -2009 255 -1941 289
rect -1851 255 -1783 289
rect -1693 255 -1625 289
rect -1535 255 -1467 289
rect -1377 255 -1309 289
rect -1219 255 -1151 289
rect -1061 255 -993 289
rect -903 255 -835 289
rect -745 255 -677 289
rect -587 255 -519 289
rect -429 255 -361 289
rect -271 255 -203 289
rect -113 255 -45 289
rect 45 255 113 289
rect 203 255 271 289
rect 361 255 429 289
rect 519 255 587 289
rect 677 255 745 289
rect 835 255 903 289
rect 993 255 1061 289
rect 1151 255 1219 289
rect 1309 255 1377 289
rect 1467 255 1535 289
rect 1625 255 1693 289
rect 1783 255 1851 289
rect 1941 255 2009 289
rect 2099 255 2167 289
rect 2257 255 2325 289
rect 2415 255 2483 289
rect 2573 255 2641 289
rect 2731 255 2799 289
rect 2889 255 2957 289
rect 3047 255 3115 289
rect 3205 255 3273 289
rect 3363 255 3431 289
rect 3521 255 3589 289
rect 3679 255 3747 289
rect 3837 255 3905 289
rect 3995 255 4063 289
rect 4153 255 4221 289
rect 4311 255 4379 289
rect -4379 147 -4311 181
rect -4221 147 -4153 181
rect -4063 147 -3995 181
rect -3905 147 -3837 181
rect -3747 147 -3679 181
rect -3589 147 -3521 181
rect -3431 147 -3363 181
rect -3273 147 -3205 181
rect -3115 147 -3047 181
rect -2957 147 -2889 181
rect -2799 147 -2731 181
rect -2641 147 -2573 181
rect -2483 147 -2415 181
rect -2325 147 -2257 181
rect -2167 147 -2099 181
rect -2009 147 -1941 181
rect -1851 147 -1783 181
rect -1693 147 -1625 181
rect -1535 147 -1467 181
rect -1377 147 -1309 181
rect -1219 147 -1151 181
rect -1061 147 -993 181
rect -903 147 -835 181
rect -745 147 -677 181
rect -587 147 -519 181
rect -429 147 -361 181
rect -271 147 -203 181
rect -113 147 -45 181
rect 45 147 113 181
rect 203 147 271 181
rect 361 147 429 181
rect 519 147 587 181
rect 677 147 745 181
rect 835 147 903 181
rect 993 147 1061 181
rect 1151 147 1219 181
rect 1309 147 1377 181
rect 1467 147 1535 181
rect 1625 147 1693 181
rect 1783 147 1851 181
rect 1941 147 2009 181
rect 2099 147 2167 181
rect 2257 147 2325 181
rect 2415 147 2483 181
rect 2573 147 2641 181
rect 2731 147 2799 181
rect 2889 147 2957 181
rect 3047 147 3115 181
rect 3205 147 3273 181
rect 3363 147 3431 181
rect 3521 147 3589 181
rect 3679 147 3747 181
rect 3837 147 3905 181
rect 3995 147 4063 181
rect 4153 147 4221 181
rect 4311 147 4379 181
rect -4379 -181 -4311 -147
rect -4221 -181 -4153 -147
rect -4063 -181 -3995 -147
rect -3905 -181 -3837 -147
rect -3747 -181 -3679 -147
rect -3589 -181 -3521 -147
rect -3431 -181 -3363 -147
rect -3273 -181 -3205 -147
rect -3115 -181 -3047 -147
rect -2957 -181 -2889 -147
rect -2799 -181 -2731 -147
rect -2641 -181 -2573 -147
rect -2483 -181 -2415 -147
rect -2325 -181 -2257 -147
rect -2167 -181 -2099 -147
rect -2009 -181 -1941 -147
rect -1851 -181 -1783 -147
rect -1693 -181 -1625 -147
rect -1535 -181 -1467 -147
rect -1377 -181 -1309 -147
rect -1219 -181 -1151 -147
rect -1061 -181 -993 -147
rect -903 -181 -835 -147
rect -745 -181 -677 -147
rect -587 -181 -519 -147
rect -429 -181 -361 -147
rect -271 -181 -203 -147
rect -113 -181 -45 -147
rect 45 -181 113 -147
rect 203 -181 271 -147
rect 361 -181 429 -147
rect 519 -181 587 -147
rect 677 -181 745 -147
rect 835 -181 903 -147
rect 993 -181 1061 -147
rect 1151 -181 1219 -147
rect 1309 -181 1377 -147
rect 1467 -181 1535 -147
rect 1625 -181 1693 -147
rect 1783 -181 1851 -147
rect 1941 -181 2009 -147
rect 2099 -181 2167 -147
rect 2257 -181 2325 -147
rect 2415 -181 2483 -147
rect 2573 -181 2641 -147
rect 2731 -181 2799 -147
rect 2889 -181 2957 -147
rect 3047 -181 3115 -147
rect 3205 -181 3273 -147
rect 3363 -181 3431 -147
rect 3521 -181 3589 -147
rect 3679 -181 3747 -147
rect 3837 -181 3905 -147
rect 3995 -181 4063 -147
rect 4153 -181 4221 -147
rect 4311 -181 4379 -147
rect -4379 -289 -4311 -255
rect -4221 -289 -4153 -255
rect -4063 -289 -3995 -255
rect -3905 -289 -3837 -255
rect -3747 -289 -3679 -255
rect -3589 -289 -3521 -255
rect -3431 -289 -3363 -255
rect -3273 -289 -3205 -255
rect -3115 -289 -3047 -255
rect -2957 -289 -2889 -255
rect -2799 -289 -2731 -255
rect -2641 -289 -2573 -255
rect -2483 -289 -2415 -255
rect -2325 -289 -2257 -255
rect -2167 -289 -2099 -255
rect -2009 -289 -1941 -255
rect -1851 -289 -1783 -255
rect -1693 -289 -1625 -255
rect -1535 -289 -1467 -255
rect -1377 -289 -1309 -255
rect -1219 -289 -1151 -255
rect -1061 -289 -993 -255
rect -903 -289 -835 -255
rect -745 -289 -677 -255
rect -587 -289 -519 -255
rect -429 -289 -361 -255
rect -271 -289 -203 -255
rect -113 -289 -45 -255
rect 45 -289 113 -255
rect 203 -289 271 -255
rect 361 -289 429 -255
rect 519 -289 587 -255
rect 677 -289 745 -255
rect 835 -289 903 -255
rect 993 -289 1061 -255
rect 1151 -289 1219 -255
rect 1309 -289 1377 -255
rect 1467 -289 1535 -255
rect 1625 -289 1693 -255
rect 1783 -289 1851 -255
rect 1941 -289 2009 -255
rect 2099 -289 2167 -255
rect 2257 -289 2325 -255
rect 2415 -289 2483 -255
rect 2573 -289 2641 -255
rect 2731 -289 2799 -255
rect 2889 -289 2957 -255
rect 3047 -289 3115 -255
rect 3205 -289 3273 -255
rect 3363 -289 3431 -255
rect 3521 -289 3589 -255
rect 3679 -289 3747 -255
rect 3837 -289 3905 -255
rect 3995 -289 4063 -255
rect 4153 -289 4221 -255
rect 4311 -289 4379 -255
rect -4379 -617 -4311 -583
rect -4221 -617 -4153 -583
rect -4063 -617 -3995 -583
rect -3905 -617 -3837 -583
rect -3747 -617 -3679 -583
rect -3589 -617 -3521 -583
rect -3431 -617 -3363 -583
rect -3273 -617 -3205 -583
rect -3115 -617 -3047 -583
rect -2957 -617 -2889 -583
rect -2799 -617 -2731 -583
rect -2641 -617 -2573 -583
rect -2483 -617 -2415 -583
rect -2325 -617 -2257 -583
rect -2167 -617 -2099 -583
rect -2009 -617 -1941 -583
rect -1851 -617 -1783 -583
rect -1693 -617 -1625 -583
rect -1535 -617 -1467 -583
rect -1377 -617 -1309 -583
rect -1219 -617 -1151 -583
rect -1061 -617 -993 -583
rect -903 -617 -835 -583
rect -745 -617 -677 -583
rect -587 -617 -519 -583
rect -429 -617 -361 -583
rect -271 -617 -203 -583
rect -113 -617 -45 -583
rect 45 -617 113 -583
rect 203 -617 271 -583
rect 361 -617 429 -583
rect 519 -617 587 -583
rect 677 -617 745 -583
rect 835 -617 903 -583
rect 993 -617 1061 -583
rect 1151 -617 1219 -583
rect 1309 -617 1377 -583
rect 1467 -617 1535 -583
rect 1625 -617 1693 -583
rect 1783 -617 1851 -583
rect 1941 -617 2009 -583
rect 2099 -617 2167 -583
rect 2257 -617 2325 -583
rect 2415 -617 2483 -583
rect 2573 -617 2641 -583
rect 2731 -617 2799 -583
rect 2889 -617 2957 -583
rect 3047 -617 3115 -583
rect 3205 -617 3273 -583
rect 3363 -617 3431 -583
rect 3521 -617 3589 -583
rect 3679 -617 3747 -583
rect 3837 -617 3905 -583
rect 3995 -617 4063 -583
rect 4153 -617 4221 -583
rect 4311 -617 4379 -583
rect -4379 -725 -4311 -691
rect -4221 -725 -4153 -691
rect -4063 -725 -3995 -691
rect -3905 -725 -3837 -691
rect -3747 -725 -3679 -691
rect -3589 -725 -3521 -691
rect -3431 -725 -3363 -691
rect -3273 -725 -3205 -691
rect -3115 -725 -3047 -691
rect -2957 -725 -2889 -691
rect -2799 -725 -2731 -691
rect -2641 -725 -2573 -691
rect -2483 -725 -2415 -691
rect -2325 -725 -2257 -691
rect -2167 -725 -2099 -691
rect -2009 -725 -1941 -691
rect -1851 -725 -1783 -691
rect -1693 -725 -1625 -691
rect -1535 -725 -1467 -691
rect -1377 -725 -1309 -691
rect -1219 -725 -1151 -691
rect -1061 -725 -993 -691
rect -903 -725 -835 -691
rect -745 -725 -677 -691
rect -587 -725 -519 -691
rect -429 -725 -361 -691
rect -271 -725 -203 -691
rect -113 -725 -45 -691
rect 45 -725 113 -691
rect 203 -725 271 -691
rect 361 -725 429 -691
rect 519 -725 587 -691
rect 677 -725 745 -691
rect 835 -725 903 -691
rect 993 -725 1061 -691
rect 1151 -725 1219 -691
rect 1309 -725 1377 -691
rect 1467 -725 1535 -691
rect 1625 -725 1693 -691
rect 1783 -725 1851 -691
rect 1941 -725 2009 -691
rect 2099 -725 2167 -691
rect 2257 -725 2325 -691
rect 2415 -725 2483 -691
rect 2573 -725 2641 -691
rect 2731 -725 2799 -691
rect 2889 -725 2957 -691
rect 3047 -725 3115 -691
rect 3205 -725 3273 -691
rect 3363 -725 3431 -691
rect 3521 -725 3589 -691
rect 3679 -725 3747 -691
rect 3837 -725 3905 -691
rect 3995 -725 4063 -691
rect 4153 -725 4221 -691
rect 4311 -725 4379 -691
rect -4379 -1053 -4311 -1019
rect -4221 -1053 -4153 -1019
rect -4063 -1053 -3995 -1019
rect -3905 -1053 -3837 -1019
rect -3747 -1053 -3679 -1019
rect -3589 -1053 -3521 -1019
rect -3431 -1053 -3363 -1019
rect -3273 -1053 -3205 -1019
rect -3115 -1053 -3047 -1019
rect -2957 -1053 -2889 -1019
rect -2799 -1053 -2731 -1019
rect -2641 -1053 -2573 -1019
rect -2483 -1053 -2415 -1019
rect -2325 -1053 -2257 -1019
rect -2167 -1053 -2099 -1019
rect -2009 -1053 -1941 -1019
rect -1851 -1053 -1783 -1019
rect -1693 -1053 -1625 -1019
rect -1535 -1053 -1467 -1019
rect -1377 -1053 -1309 -1019
rect -1219 -1053 -1151 -1019
rect -1061 -1053 -993 -1019
rect -903 -1053 -835 -1019
rect -745 -1053 -677 -1019
rect -587 -1053 -519 -1019
rect -429 -1053 -361 -1019
rect -271 -1053 -203 -1019
rect -113 -1053 -45 -1019
rect 45 -1053 113 -1019
rect 203 -1053 271 -1019
rect 361 -1053 429 -1019
rect 519 -1053 587 -1019
rect 677 -1053 745 -1019
rect 835 -1053 903 -1019
rect 993 -1053 1061 -1019
rect 1151 -1053 1219 -1019
rect 1309 -1053 1377 -1019
rect 1467 -1053 1535 -1019
rect 1625 -1053 1693 -1019
rect 1783 -1053 1851 -1019
rect 1941 -1053 2009 -1019
rect 2099 -1053 2167 -1019
rect 2257 -1053 2325 -1019
rect 2415 -1053 2483 -1019
rect 2573 -1053 2641 -1019
rect 2731 -1053 2799 -1019
rect 2889 -1053 2957 -1019
rect 3047 -1053 3115 -1019
rect 3205 -1053 3273 -1019
rect 3363 -1053 3431 -1019
rect 3521 -1053 3589 -1019
rect 3679 -1053 3747 -1019
rect 3837 -1053 3905 -1019
rect 3995 -1053 4063 -1019
rect 4153 -1053 4221 -1019
rect 4311 -1053 4379 -1019
<< locali >>
rect -4575 1157 -4479 1191
rect 4479 1157 4575 1191
rect -4575 1095 -4541 1157
rect 4541 1095 4575 1157
rect -4395 1019 -4379 1053
rect -4311 1019 -4295 1053
rect -4237 1019 -4221 1053
rect -4153 1019 -4137 1053
rect -4079 1019 -4063 1053
rect -3995 1019 -3979 1053
rect -3921 1019 -3905 1053
rect -3837 1019 -3821 1053
rect -3763 1019 -3747 1053
rect -3679 1019 -3663 1053
rect -3605 1019 -3589 1053
rect -3521 1019 -3505 1053
rect -3447 1019 -3431 1053
rect -3363 1019 -3347 1053
rect -3289 1019 -3273 1053
rect -3205 1019 -3189 1053
rect -3131 1019 -3115 1053
rect -3047 1019 -3031 1053
rect -2973 1019 -2957 1053
rect -2889 1019 -2873 1053
rect -2815 1019 -2799 1053
rect -2731 1019 -2715 1053
rect -2657 1019 -2641 1053
rect -2573 1019 -2557 1053
rect -2499 1019 -2483 1053
rect -2415 1019 -2399 1053
rect -2341 1019 -2325 1053
rect -2257 1019 -2241 1053
rect -2183 1019 -2167 1053
rect -2099 1019 -2083 1053
rect -2025 1019 -2009 1053
rect -1941 1019 -1925 1053
rect -1867 1019 -1851 1053
rect -1783 1019 -1767 1053
rect -1709 1019 -1693 1053
rect -1625 1019 -1609 1053
rect -1551 1019 -1535 1053
rect -1467 1019 -1451 1053
rect -1393 1019 -1377 1053
rect -1309 1019 -1293 1053
rect -1235 1019 -1219 1053
rect -1151 1019 -1135 1053
rect -1077 1019 -1061 1053
rect -993 1019 -977 1053
rect -919 1019 -903 1053
rect -835 1019 -819 1053
rect -761 1019 -745 1053
rect -677 1019 -661 1053
rect -603 1019 -587 1053
rect -519 1019 -503 1053
rect -445 1019 -429 1053
rect -361 1019 -345 1053
rect -287 1019 -271 1053
rect -203 1019 -187 1053
rect -129 1019 -113 1053
rect -45 1019 -29 1053
rect 29 1019 45 1053
rect 113 1019 129 1053
rect 187 1019 203 1053
rect 271 1019 287 1053
rect 345 1019 361 1053
rect 429 1019 445 1053
rect 503 1019 519 1053
rect 587 1019 603 1053
rect 661 1019 677 1053
rect 745 1019 761 1053
rect 819 1019 835 1053
rect 903 1019 919 1053
rect 977 1019 993 1053
rect 1061 1019 1077 1053
rect 1135 1019 1151 1053
rect 1219 1019 1235 1053
rect 1293 1019 1309 1053
rect 1377 1019 1393 1053
rect 1451 1019 1467 1053
rect 1535 1019 1551 1053
rect 1609 1019 1625 1053
rect 1693 1019 1709 1053
rect 1767 1019 1783 1053
rect 1851 1019 1867 1053
rect 1925 1019 1941 1053
rect 2009 1019 2025 1053
rect 2083 1019 2099 1053
rect 2167 1019 2183 1053
rect 2241 1019 2257 1053
rect 2325 1019 2341 1053
rect 2399 1019 2415 1053
rect 2483 1019 2499 1053
rect 2557 1019 2573 1053
rect 2641 1019 2657 1053
rect 2715 1019 2731 1053
rect 2799 1019 2815 1053
rect 2873 1019 2889 1053
rect 2957 1019 2973 1053
rect 3031 1019 3047 1053
rect 3115 1019 3131 1053
rect 3189 1019 3205 1053
rect 3273 1019 3289 1053
rect 3347 1019 3363 1053
rect 3431 1019 3447 1053
rect 3505 1019 3521 1053
rect 3589 1019 3605 1053
rect 3663 1019 3679 1053
rect 3747 1019 3763 1053
rect 3821 1019 3837 1053
rect 3905 1019 3921 1053
rect 3979 1019 3995 1053
rect 4063 1019 4079 1053
rect 4137 1019 4153 1053
rect 4221 1019 4237 1053
rect 4295 1019 4311 1053
rect 4379 1019 4395 1053
rect -4441 960 -4407 976
rect -4441 768 -4407 784
rect -4283 960 -4249 976
rect -4283 768 -4249 784
rect -4125 960 -4091 976
rect -4125 768 -4091 784
rect -3967 960 -3933 976
rect -3967 768 -3933 784
rect -3809 960 -3775 976
rect -3809 768 -3775 784
rect -3651 960 -3617 976
rect -3651 768 -3617 784
rect -3493 960 -3459 976
rect -3493 768 -3459 784
rect -3335 960 -3301 976
rect -3335 768 -3301 784
rect -3177 960 -3143 976
rect -3177 768 -3143 784
rect -3019 960 -2985 976
rect -3019 768 -2985 784
rect -2861 960 -2827 976
rect -2861 768 -2827 784
rect -2703 960 -2669 976
rect -2703 768 -2669 784
rect -2545 960 -2511 976
rect -2545 768 -2511 784
rect -2387 960 -2353 976
rect -2387 768 -2353 784
rect -2229 960 -2195 976
rect -2229 768 -2195 784
rect -2071 960 -2037 976
rect -2071 768 -2037 784
rect -1913 960 -1879 976
rect -1913 768 -1879 784
rect -1755 960 -1721 976
rect -1755 768 -1721 784
rect -1597 960 -1563 976
rect -1597 768 -1563 784
rect -1439 960 -1405 976
rect -1439 768 -1405 784
rect -1281 960 -1247 976
rect -1281 768 -1247 784
rect -1123 960 -1089 976
rect -1123 768 -1089 784
rect -965 960 -931 976
rect -965 768 -931 784
rect -807 960 -773 976
rect -807 768 -773 784
rect -649 960 -615 976
rect -649 768 -615 784
rect -491 960 -457 976
rect -491 768 -457 784
rect -333 960 -299 976
rect -333 768 -299 784
rect -175 960 -141 976
rect -175 768 -141 784
rect -17 960 17 976
rect -17 768 17 784
rect 141 960 175 976
rect 141 768 175 784
rect 299 960 333 976
rect 299 768 333 784
rect 457 960 491 976
rect 457 768 491 784
rect 615 960 649 976
rect 615 768 649 784
rect 773 960 807 976
rect 773 768 807 784
rect 931 960 965 976
rect 931 768 965 784
rect 1089 960 1123 976
rect 1089 768 1123 784
rect 1247 960 1281 976
rect 1247 768 1281 784
rect 1405 960 1439 976
rect 1405 768 1439 784
rect 1563 960 1597 976
rect 1563 768 1597 784
rect 1721 960 1755 976
rect 1721 768 1755 784
rect 1879 960 1913 976
rect 1879 768 1913 784
rect 2037 960 2071 976
rect 2037 768 2071 784
rect 2195 960 2229 976
rect 2195 768 2229 784
rect 2353 960 2387 976
rect 2353 768 2387 784
rect 2511 960 2545 976
rect 2511 768 2545 784
rect 2669 960 2703 976
rect 2669 768 2703 784
rect 2827 960 2861 976
rect 2827 768 2861 784
rect 2985 960 3019 976
rect 2985 768 3019 784
rect 3143 960 3177 976
rect 3143 768 3177 784
rect 3301 960 3335 976
rect 3301 768 3335 784
rect 3459 960 3493 976
rect 3459 768 3493 784
rect 3617 960 3651 976
rect 3617 768 3651 784
rect 3775 960 3809 976
rect 3775 768 3809 784
rect 3933 960 3967 976
rect 3933 768 3967 784
rect 4091 960 4125 976
rect 4091 768 4125 784
rect 4249 960 4283 976
rect 4249 768 4283 784
rect 4407 960 4441 976
rect 4407 768 4441 784
rect -4395 691 -4379 725
rect -4311 691 -4295 725
rect -4237 691 -4221 725
rect -4153 691 -4137 725
rect -4079 691 -4063 725
rect -3995 691 -3979 725
rect -3921 691 -3905 725
rect -3837 691 -3821 725
rect -3763 691 -3747 725
rect -3679 691 -3663 725
rect -3605 691 -3589 725
rect -3521 691 -3505 725
rect -3447 691 -3431 725
rect -3363 691 -3347 725
rect -3289 691 -3273 725
rect -3205 691 -3189 725
rect -3131 691 -3115 725
rect -3047 691 -3031 725
rect -2973 691 -2957 725
rect -2889 691 -2873 725
rect -2815 691 -2799 725
rect -2731 691 -2715 725
rect -2657 691 -2641 725
rect -2573 691 -2557 725
rect -2499 691 -2483 725
rect -2415 691 -2399 725
rect -2341 691 -2325 725
rect -2257 691 -2241 725
rect -2183 691 -2167 725
rect -2099 691 -2083 725
rect -2025 691 -2009 725
rect -1941 691 -1925 725
rect -1867 691 -1851 725
rect -1783 691 -1767 725
rect -1709 691 -1693 725
rect -1625 691 -1609 725
rect -1551 691 -1535 725
rect -1467 691 -1451 725
rect -1393 691 -1377 725
rect -1309 691 -1293 725
rect -1235 691 -1219 725
rect -1151 691 -1135 725
rect -1077 691 -1061 725
rect -993 691 -977 725
rect -919 691 -903 725
rect -835 691 -819 725
rect -761 691 -745 725
rect -677 691 -661 725
rect -603 691 -587 725
rect -519 691 -503 725
rect -445 691 -429 725
rect -361 691 -345 725
rect -287 691 -271 725
rect -203 691 -187 725
rect -129 691 -113 725
rect -45 691 -29 725
rect 29 691 45 725
rect 113 691 129 725
rect 187 691 203 725
rect 271 691 287 725
rect 345 691 361 725
rect 429 691 445 725
rect 503 691 519 725
rect 587 691 603 725
rect 661 691 677 725
rect 745 691 761 725
rect 819 691 835 725
rect 903 691 919 725
rect 977 691 993 725
rect 1061 691 1077 725
rect 1135 691 1151 725
rect 1219 691 1235 725
rect 1293 691 1309 725
rect 1377 691 1393 725
rect 1451 691 1467 725
rect 1535 691 1551 725
rect 1609 691 1625 725
rect 1693 691 1709 725
rect 1767 691 1783 725
rect 1851 691 1867 725
rect 1925 691 1941 725
rect 2009 691 2025 725
rect 2083 691 2099 725
rect 2167 691 2183 725
rect 2241 691 2257 725
rect 2325 691 2341 725
rect 2399 691 2415 725
rect 2483 691 2499 725
rect 2557 691 2573 725
rect 2641 691 2657 725
rect 2715 691 2731 725
rect 2799 691 2815 725
rect 2873 691 2889 725
rect 2957 691 2973 725
rect 3031 691 3047 725
rect 3115 691 3131 725
rect 3189 691 3205 725
rect 3273 691 3289 725
rect 3347 691 3363 725
rect 3431 691 3447 725
rect 3505 691 3521 725
rect 3589 691 3605 725
rect 3663 691 3679 725
rect 3747 691 3763 725
rect 3821 691 3837 725
rect 3905 691 3921 725
rect 3979 691 3995 725
rect 4063 691 4079 725
rect 4137 691 4153 725
rect 4221 691 4237 725
rect 4295 691 4311 725
rect 4379 691 4395 725
rect -4395 583 -4379 617
rect -4311 583 -4295 617
rect -4237 583 -4221 617
rect -4153 583 -4137 617
rect -4079 583 -4063 617
rect -3995 583 -3979 617
rect -3921 583 -3905 617
rect -3837 583 -3821 617
rect -3763 583 -3747 617
rect -3679 583 -3663 617
rect -3605 583 -3589 617
rect -3521 583 -3505 617
rect -3447 583 -3431 617
rect -3363 583 -3347 617
rect -3289 583 -3273 617
rect -3205 583 -3189 617
rect -3131 583 -3115 617
rect -3047 583 -3031 617
rect -2973 583 -2957 617
rect -2889 583 -2873 617
rect -2815 583 -2799 617
rect -2731 583 -2715 617
rect -2657 583 -2641 617
rect -2573 583 -2557 617
rect -2499 583 -2483 617
rect -2415 583 -2399 617
rect -2341 583 -2325 617
rect -2257 583 -2241 617
rect -2183 583 -2167 617
rect -2099 583 -2083 617
rect -2025 583 -2009 617
rect -1941 583 -1925 617
rect -1867 583 -1851 617
rect -1783 583 -1767 617
rect -1709 583 -1693 617
rect -1625 583 -1609 617
rect -1551 583 -1535 617
rect -1467 583 -1451 617
rect -1393 583 -1377 617
rect -1309 583 -1293 617
rect -1235 583 -1219 617
rect -1151 583 -1135 617
rect -1077 583 -1061 617
rect -993 583 -977 617
rect -919 583 -903 617
rect -835 583 -819 617
rect -761 583 -745 617
rect -677 583 -661 617
rect -603 583 -587 617
rect -519 583 -503 617
rect -445 583 -429 617
rect -361 583 -345 617
rect -287 583 -271 617
rect -203 583 -187 617
rect -129 583 -113 617
rect -45 583 -29 617
rect 29 583 45 617
rect 113 583 129 617
rect 187 583 203 617
rect 271 583 287 617
rect 345 583 361 617
rect 429 583 445 617
rect 503 583 519 617
rect 587 583 603 617
rect 661 583 677 617
rect 745 583 761 617
rect 819 583 835 617
rect 903 583 919 617
rect 977 583 993 617
rect 1061 583 1077 617
rect 1135 583 1151 617
rect 1219 583 1235 617
rect 1293 583 1309 617
rect 1377 583 1393 617
rect 1451 583 1467 617
rect 1535 583 1551 617
rect 1609 583 1625 617
rect 1693 583 1709 617
rect 1767 583 1783 617
rect 1851 583 1867 617
rect 1925 583 1941 617
rect 2009 583 2025 617
rect 2083 583 2099 617
rect 2167 583 2183 617
rect 2241 583 2257 617
rect 2325 583 2341 617
rect 2399 583 2415 617
rect 2483 583 2499 617
rect 2557 583 2573 617
rect 2641 583 2657 617
rect 2715 583 2731 617
rect 2799 583 2815 617
rect 2873 583 2889 617
rect 2957 583 2973 617
rect 3031 583 3047 617
rect 3115 583 3131 617
rect 3189 583 3205 617
rect 3273 583 3289 617
rect 3347 583 3363 617
rect 3431 583 3447 617
rect 3505 583 3521 617
rect 3589 583 3605 617
rect 3663 583 3679 617
rect 3747 583 3763 617
rect 3821 583 3837 617
rect 3905 583 3921 617
rect 3979 583 3995 617
rect 4063 583 4079 617
rect 4137 583 4153 617
rect 4221 583 4237 617
rect 4295 583 4311 617
rect 4379 583 4395 617
rect -4441 524 -4407 540
rect -4441 332 -4407 348
rect -4283 524 -4249 540
rect -4283 332 -4249 348
rect -4125 524 -4091 540
rect -4125 332 -4091 348
rect -3967 524 -3933 540
rect -3967 332 -3933 348
rect -3809 524 -3775 540
rect -3809 332 -3775 348
rect -3651 524 -3617 540
rect -3651 332 -3617 348
rect -3493 524 -3459 540
rect -3493 332 -3459 348
rect -3335 524 -3301 540
rect -3335 332 -3301 348
rect -3177 524 -3143 540
rect -3177 332 -3143 348
rect -3019 524 -2985 540
rect -3019 332 -2985 348
rect -2861 524 -2827 540
rect -2861 332 -2827 348
rect -2703 524 -2669 540
rect -2703 332 -2669 348
rect -2545 524 -2511 540
rect -2545 332 -2511 348
rect -2387 524 -2353 540
rect -2387 332 -2353 348
rect -2229 524 -2195 540
rect -2229 332 -2195 348
rect -2071 524 -2037 540
rect -2071 332 -2037 348
rect -1913 524 -1879 540
rect -1913 332 -1879 348
rect -1755 524 -1721 540
rect -1755 332 -1721 348
rect -1597 524 -1563 540
rect -1597 332 -1563 348
rect -1439 524 -1405 540
rect -1439 332 -1405 348
rect -1281 524 -1247 540
rect -1281 332 -1247 348
rect -1123 524 -1089 540
rect -1123 332 -1089 348
rect -965 524 -931 540
rect -965 332 -931 348
rect -807 524 -773 540
rect -807 332 -773 348
rect -649 524 -615 540
rect -649 332 -615 348
rect -491 524 -457 540
rect -491 332 -457 348
rect -333 524 -299 540
rect -333 332 -299 348
rect -175 524 -141 540
rect -175 332 -141 348
rect -17 524 17 540
rect -17 332 17 348
rect 141 524 175 540
rect 141 332 175 348
rect 299 524 333 540
rect 299 332 333 348
rect 457 524 491 540
rect 457 332 491 348
rect 615 524 649 540
rect 615 332 649 348
rect 773 524 807 540
rect 773 332 807 348
rect 931 524 965 540
rect 931 332 965 348
rect 1089 524 1123 540
rect 1089 332 1123 348
rect 1247 524 1281 540
rect 1247 332 1281 348
rect 1405 524 1439 540
rect 1405 332 1439 348
rect 1563 524 1597 540
rect 1563 332 1597 348
rect 1721 524 1755 540
rect 1721 332 1755 348
rect 1879 524 1913 540
rect 1879 332 1913 348
rect 2037 524 2071 540
rect 2037 332 2071 348
rect 2195 524 2229 540
rect 2195 332 2229 348
rect 2353 524 2387 540
rect 2353 332 2387 348
rect 2511 524 2545 540
rect 2511 332 2545 348
rect 2669 524 2703 540
rect 2669 332 2703 348
rect 2827 524 2861 540
rect 2827 332 2861 348
rect 2985 524 3019 540
rect 2985 332 3019 348
rect 3143 524 3177 540
rect 3143 332 3177 348
rect 3301 524 3335 540
rect 3301 332 3335 348
rect 3459 524 3493 540
rect 3459 332 3493 348
rect 3617 524 3651 540
rect 3617 332 3651 348
rect 3775 524 3809 540
rect 3775 332 3809 348
rect 3933 524 3967 540
rect 3933 332 3967 348
rect 4091 524 4125 540
rect 4091 332 4125 348
rect 4249 524 4283 540
rect 4249 332 4283 348
rect 4407 524 4441 540
rect 4407 332 4441 348
rect -4395 255 -4379 289
rect -4311 255 -4295 289
rect -4237 255 -4221 289
rect -4153 255 -4137 289
rect -4079 255 -4063 289
rect -3995 255 -3979 289
rect -3921 255 -3905 289
rect -3837 255 -3821 289
rect -3763 255 -3747 289
rect -3679 255 -3663 289
rect -3605 255 -3589 289
rect -3521 255 -3505 289
rect -3447 255 -3431 289
rect -3363 255 -3347 289
rect -3289 255 -3273 289
rect -3205 255 -3189 289
rect -3131 255 -3115 289
rect -3047 255 -3031 289
rect -2973 255 -2957 289
rect -2889 255 -2873 289
rect -2815 255 -2799 289
rect -2731 255 -2715 289
rect -2657 255 -2641 289
rect -2573 255 -2557 289
rect -2499 255 -2483 289
rect -2415 255 -2399 289
rect -2341 255 -2325 289
rect -2257 255 -2241 289
rect -2183 255 -2167 289
rect -2099 255 -2083 289
rect -2025 255 -2009 289
rect -1941 255 -1925 289
rect -1867 255 -1851 289
rect -1783 255 -1767 289
rect -1709 255 -1693 289
rect -1625 255 -1609 289
rect -1551 255 -1535 289
rect -1467 255 -1451 289
rect -1393 255 -1377 289
rect -1309 255 -1293 289
rect -1235 255 -1219 289
rect -1151 255 -1135 289
rect -1077 255 -1061 289
rect -993 255 -977 289
rect -919 255 -903 289
rect -835 255 -819 289
rect -761 255 -745 289
rect -677 255 -661 289
rect -603 255 -587 289
rect -519 255 -503 289
rect -445 255 -429 289
rect -361 255 -345 289
rect -287 255 -271 289
rect -203 255 -187 289
rect -129 255 -113 289
rect -45 255 -29 289
rect 29 255 45 289
rect 113 255 129 289
rect 187 255 203 289
rect 271 255 287 289
rect 345 255 361 289
rect 429 255 445 289
rect 503 255 519 289
rect 587 255 603 289
rect 661 255 677 289
rect 745 255 761 289
rect 819 255 835 289
rect 903 255 919 289
rect 977 255 993 289
rect 1061 255 1077 289
rect 1135 255 1151 289
rect 1219 255 1235 289
rect 1293 255 1309 289
rect 1377 255 1393 289
rect 1451 255 1467 289
rect 1535 255 1551 289
rect 1609 255 1625 289
rect 1693 255 1709 289
rect 1767 255 1783 289
rect 1851 255 1867 289
rect 1925 255 1941 289
rect 2009 255 2025 289
rect 2083 255 2099 289
rect 2167 255 2183 289
rect 2241 255 2257 289
rect 2325 255 2341 289
rect 2399 255 2415 289
rect 2483 255 2499 289
rect 2557 255 2573 289
rect 2641 255 2657 289
rect 2715 255 2731 289
rect 2799 255 2815 289
rect 2873 255 2889 289
rect 2957 255 2973 289
rect 3031 255 3047 289
rect 3115 255 3131 289
rect 3189 255 3205 289
rect 3273 255 3289 289
rect 3347 255 3363 289
rect 3431 255 3447 289
rect 3505 255 3521 289
rect 3589 255 3605 289
rect 3663 255 3679 289
rect 3747 255 3763 289
rect 3821 255 3837 289
rect 3905 255 3921 289
rect 3979 255 3995 289
rect 4063 255 4079 289
rect 4137 255 4153 289
rect 4221 255 4237 289
rect 4295 255 4311 289
rect 4379 255 4395 289
rect -4395 147 -4379 181
rect -4311 147 -4295 181
rect -4237 147 -4221 181
rect -4153 147 -4137 181
rect -4079 147 -4063 181
rect -3995 147 -3979 181
rect -3921 147 -3905 181
rect -3837 147 -3821 181
rect -3763 147 -3747 181
rect -3679 147 -3663 181
rect -3605 147 -3589 181
rect -3521 147 -3505 181
rect -3447 147 -3431 181
rect -3363 147 -3347 181
rect -3289 147 -3273 181
rect -3205 147 -3189 181
rect -3131 147 -3115 181
rect -3047 147 -3031 181
rect -2973 147 -2957 181
rect -2889 147 -2873 181
rect -2815 147 -2799 181
rect -2731 147 -2715 181
rect -2657 147 -2641 181
rect -2573 147 -2557 181
rect -2499 147 -2483 181
rect -2415 147 -2399 181
rect -2341 147 -2325 181
rect -2257 147 -2241 181
rect -2183 147 -2167 181
rect -2099 147 -2083 181
rect -2025 147 -2009 181
rect -1941 147 -1925 181
rect -1867 147 -1851 181
rect -1783 147 -1767 181
rect -1709 147 -1693 181
rect -1625 147 -1609 181
rect -1551 147 -1535 181
rect -1467 147 -1451 181
rect -1393 147 -1377 181
rect -1309 147 -1293 181
rect -1235 147 -1219 181
rect -1151 147 -1135 181
rect -1077 147 -1061 181
rect -993 147 -977 181
rect -919 147 -903 181
rect -835 147 -819 181
rect -761 147 -745 181
rect -677 147 -661 181
rect -603 147 -587 181
rect -519 147 -503 181
rect -445 147 -429 181
rect -361 147 -345 181
rect -287 147 -271 181
rect -203 147 -187 181
rect -129 147 -113 181
rect -45 147 -29 181
rect 29 147 45 181
rect 113 147 129 181
rect 187 147 203 181
rect 271 147 287 181
rect 345 147 361 181
rect 429 147 445 181
rect 503 147 519 181
rect 587 147 603 181
rect 661 147 677 181
rect 745 147 761 181
rect 819 147 835 181
rect 903 147 919 181
rect 977 147 993 181
rect 1061 147 1077 181
rect 1135 147 1151 181
rect 1219 147 1235 181
rect 1293 147 1309 181
rect 1377 147 1393 181
rect 1451 147 1467 181
rect 1535 147 1551 181
rect 1609 147 1625 181
rect 1693 147 1709 181
rect 1767 147 1783 181
rect 1851 147 1867 181
rect 1925 147 1941 181
rect 2009 147 2025 181
rect 2083 147 2099 181
rect 2167 147 2183 181
rect 2241 147 2257 181
rect 2325 147 2341 181
rect 2399 147 2415 181
rect 2483 147 2499 181
rect 2557 147 2573 181
rect 2641 147 2657 181
rect 2715 147 2731 181
rect 2799 147 2815 181
rect 2873 147 2889 181
rect 2957 147 2973 181
rect 3031 147 3047 181
rect 3115 147 3131 181
rect 3189 147 3205 181
rect 3273 147 3289 181
rect 3347 147 3363 181
rect 3431 147 3447 181
rect 3505 147 3521 181
rect 3589 147 3605 181
rect 3663 147 3679 181
rect 3747 147 3763 181
rect 3821 147 3837 181
rect 3905 147 3921 181
rect 3979 147 3995 181
rect 4063 147 4079 181
rect 4137 147 4153 181
rect 4221 147 4237 181
rect 4295 147 4311 181
rect 4379 147 4395 181
rect -4441 88 -4407 104
rect -4441 -104 -4407 -88
rect -4283 88 -4249 104
rect -4283 -104 -4249 -88
rect -4125 88 -4091 104
rect -4125 -104 -4091 -88
rect -3967 88 -3933 104
rect -3967 -104 -3933 -88
rect -3809 88 -3775 104
rect -3809 -104 -3775 -88
rect -3651 88 -3617 104
rect -3651 -104 -3617 -88
rect -3493 88 -3459 104
rect -3493 -104 -3459 -88
rect -3335 88 -3301 104
rect -3335 -104 -3301 -88
rect -3177 88 -3143 104
rect -3177 -104 -3143 -88
rect -3019 88 -2985 104
rect -3019 -104 -2985 -88
rect -2861 88 -2827 104
rect -2861 -104 -2827 -88
rect -2703 88 -2669 104
rect -2703 -104 -2669 -88
rect -2545 88 -2511 104
rect -2545 -104 -2511 -88
rect -2387 88 -2353 104
rect -2387 -104 -2353 -88
rect -2229 88 -2195 104
rect -2229 -104 -2195 -88
rect -2071 88 -2037 104
rect -2071 -104 -2037 -88
rect -1913 88 -1879 104
rect -1913 -104 -1879 -88
rect -1755 88 -1721 104
rect -1755 -104 -1721 -88
rect -1597 88 -1563 104
rect -1597 -104 -1563 -88
rect -1439 88 -1405 104
rect -1439 -104 -1405 -88
rect -1281 88 -1247 104
rect -1281 -104 -1247 -88
rect -1123 88 -1089 104
rect -1123 -104 -1089 -88
rect -965 88 -931 104
rect -965 -104 -931 -88
rect -807 88 -773 104
rect -807 -104 -773 -88
rect -649 88 -615 104
rect -649 -104 -615 -88
rect -491 88 -457 104
rect -491 -104 -457 -88
rect -333 88 -299 104
rect -333 -104 -299 -88
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect 299 88 333 104
rect 299 -104 333 -88
rect 457 88 491 104
rect 457 -104 491 -88
rect 615 88 649 104
rect 615 -104 649 -88
rect 773 88 807 104
rect 773 -104 807 -88
rect 931 88 965 104
rect 931 -104 965 -88
rect 1089 88 1123 104
rect 1089 -104 1123 -88
rect 1247 88 1281 104
rect 1247 -104 1281 -88
rect 1405 88 1439 104
rect 1405 -104 1439 -88
rect 1563 88 1597 104
rect 1563 -104 1597 -88
rect 1721 88 1755 104
rect 1721 -104 1755 -88
rect 1879 88 1913 104
rect 1879 -104 1913 -88
rect 2037 88 2071 104
rect 2037 -104 2071 -88
rect 2195 88 2229 104
rect 2195 -104 2229 -88
rect 2353 88 2387 104
rect 2353 -104 2387 -88
rect 2511 88 2545 104
rect 2511 -104 2545 -88
rect 2669 88 2703 104
rect 2669 -104 2703 -88
rect 2827 88 2861 104
rect 2827 -104 2861 -88
rect 2985 88 3019 104
rect 2985 -104 3019 -88
rect 3143 88 3177 104
rect 3143 -104 3177 -88
rect 3301 88 3335 104
rect 3301 -104 3335 -88
rect 3459 88 3493 104
rect 3459 -104 3493 -88
rect 3617 88 3651 104
rect 3617 -104 3651 -88
rect 3775 88 3809 104
rect 3775 -104 3809 -88
rect 3933 88 3967 104
rect 3933 -104 3967 -88
rect 4091 88 4125 104
rect 4091 -104 4125 -88
rect 4249 88 4283 104
rect 4249 -104 4283 -88
rect 4407 88 4441 104
rect 4407 -104 4441 -88
rect -4395 -181 -4379 -147
rect -4311 -181 -4295 -147
rect -4237 -181 -4221 -147
rect -4153 -181 -4137 -147
rect -4079 -181 -4063 -147
rect -3995 -181 -3979 -147
rect -3921 -181 -3905 -147
rect -3837 -181 -3821 -147
rect -3763 -181 -3747 -147
rect -3679 -181 -3663 -147
rect -3605 -181 -3589 -147
rect -3521 -181 -3505 -147
rect -3447 -181 -3431 -147
rect -3363 -181 -3347 -147
rect -3289 -181 -3273 -147
rect -3205 -181 -3189 -147
rect -3131 -181 -3115 -147
rect -3047 -181 -3031 -147
rect -2973 -181 -2957 -147
rect -2889 -181 -2873 -147
rect -2815 -181 -2799 -147
rect -2731 -181 -2715 -147
rect -2657 -181 -2641 -147
rect -2573 -181 -2557 -147
rect -2499 -181 -2483 -147
rect -2415 -181 -2399 -147
rect -2341 -181 -2325 -147
rect -2257 -181 -2241 -147
rect -2183 -181 -2167 -147
rect -2099 -181 -2083 -147
rect -2025 -181 -2009 -147
rect -1941 -181 -1925 -147
rect -1867 -181 -1851 -147
rect -1783 -181 -1767 -147
rect -1709 -181 -1693 -147
rect -1625 -181 -1609 -147
rect -1551 -181 -1535 -147
rect -1467 -181 -1451 -147
rect -1393 -181 -1377 -147
rect -1309 -181 -1293 -147
rect -1235 -181 -1219 -147
rect -1151 -181 -1135 -147
rect -1077 -181 -1061 -147
rect -993 -181 -977 -147
rect -919 -181 -903 -147
rect -835 -181 -819 -147
rect -761 -181 -745 -147
rect -677 -181 -661 -147
rect -603 -181 -587 -147
rect -519 -181 -503 -147
rect -445 -181 -429 -147
rect -361 -181 -345 -147
rect -287 -181 -271 -147
rect -203 -181 -187 -147
rect -129 -181 -113 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 113 -181 129 -147
rect 187 -181 203 -147
rect 271 -181 287 -147
rect 345 -181 361 -147
rect 429 -181 445 -147
rect 503 -181 519 -147
rect 587 -181 603 -147
rect 661 -181 677 -147
rect 745 -181 761 -147
rect 819 -181 835 -147
rect 903 -181 919 -147
rect 977 -181 993 -147
rect 1061 -181 1077 -147
rect 1135 -181 1151 -147
rect 1219 -181 1235 -147
rect 1293 -181 1309 -147
rect 1377 -181 1393 -147
rect 1451 -181 1467 -147
rect 1535 -181 1551 -147
rect 1609 -181 1625 -147
rect 1693 -181 1709 -147
rect 1767 -181 1783 -147
rect 1851 -181 1867 -147
rect 1925 -181 1941 -147
rect 2009 -181 2025 -147
rect 2083 -181 2099 -147
rect 2167 -181 2183 -147
rect 2241 -181 2257 -147
rect 2325 -181 2341 -147
rect 2399 -181 2415 -147
rect 2483 -181 2499 -147
rect 2557 -181 2573 -147
rect 2641 -181 2657 -147
rect 2715 -181 2731 -147
rect 2799 -181 2815 -147
rect 2873 -181 2889 -147
rect 2957 -181 2973 -147
rect 3031 -181 3047 -147
rect 3115 -181 3131 -147
rect 3189 -181 3205 -147
rect 3273 -181 3289 -147
rect 3347 -181 3363 -147
rect 3431 -181 3447 -147
rect 3505 -181 3521 -147
rect 3589 -181 3605 -147
rect 3663 -181 3679 -147
rect 3747 -181 3763 -147
rect 3821 -181 3837 -147
rect 3905 -181 3921 -147
rect 3979 -181 3995 -147
rect 4063 -181 4079 -147
rect 4137 -181 4153 -147
rect 4221 -181 4237 -147
rect 4295 -181 4311 -147
rect 4379 -181 4395 -147
rect -4395 -289 -4379 -255
rect -4311 -289 -4295 -255
rect -4237 -289 -4221 -255
rect -4153 -289 -4137 -255
rect -4079 -289 -4063 -255
rect -3995 -289 -3979 -255
rect -3921 -289 -3905 -255
rect -3837 -289 -3821 -255
rect -3763 -289 -3747 -255
rect -3679 -289 -3663 -255
rect -3605 -289 -3589 -255
rect -3521 -289 -3505 -255
rect -3447 -289 -3431 -255
rect -3363 -289 -3347 -255
rect -3289 -289 -3273 -255
rect -3205 -289 -3189 -255
rect -3131 -289 -3115 -255
rect -3047 -289 -3031 -255
rect -2973 -289 -2957 -255
rect -2889 -289 -2873 -255
rect -2815 -289 -2799 -255
rect -2731 -289 -2715 -255
rect -2657 -289 -2641 -255
rect -2573 -289 -2557 -255
rect -2499 -289 -2483 -255
rect -2415 -289 -2399 -255
rect -2341 -289 -2325 -255
rect -2257 -289 -2241 -255
rect -2183 -289 -2167 -255
rect -2099 -289 -2083 -255
rect -2025 -289 -2009 -255
rect -1941 -289 -1925 -255
rect -1867 -289 -1851 -255
rect -1783 -289 -1767 -255
rect -1709 -289 -1693 -255
rect -1625 -289 -1609 -255
rect -1551 -289 -1535 -255
rect -1467 -289 -1451 -255
rect -1393 -289 -1377 -255
rect -1309 -289 -1293 -255
rect -1235 -289 -1219 -255
rect -1151 -289 -1135 -255
rect -1077 -289 -1061 -255
rect -993 -289 -977 -255
rect -919 -289 -903 -255
rect -835 -289 -819 -255
rect -761 -289 -745 -255
rect -677 -289 -661 -255
rect -603 -289 -587 -255
rect -519 -289 -503 -255
rect -445 -289 -429 -255
rect -361 -289 -345 -255
rect -287 -289 -271 -255
rect -203 -289 -187 -255
rect -129 -289 -113 -255
rect -45 -289 -29 -255
rect 29 -289 45 -255
rect 113 -289 129 -255
rect 187 -289 203 -255
rect 271 -289 287 -255
rect 345 -289 361 -255
rect 429 -289 445 -255
rect 503 -289 519 -255
rect 587 -289 603 -255
rect 661 -289 677 -255
rect 745 -289 761 -255
rect 819 -289 835 -255
rect 903 -289 919 -255
rect 977 -289 993 -255
rect 1061 -289 1077 -255
rect 1135 -289 1151 -255
rect 1219 -289 1235 -255
rect 1293 -289 1309 -255
rect 1377 -289 1393 -255
rect 1451 -289 1467 -255
rect 1535 -289 1551 -255
rect 1609 -289 1625 -255
rect 1693 -289 1709 -255
rect 1767 -289 1783 -255
rect 1851 -289 1867 -255
rect 1925 -289 1941 -255
rect 2009 -289 2025 -255
rect 2083 -289 2099 -255
rect 2167 -289 2183 -255
rect 2241 -289 2257 -255
rect 2325 -289 2341 -255
rect 2399 -289 2415 -255
rect 2483 -289 2499 -255
rect 2557 -289 2573 -255
rect 2641 -289 2657 -255
rect 2715 -289 2731 -255
rect 2799 -289 2815 -255
rect 2873 -289 2889 -255
rect 2957 -289 2973 -255
rect 3031 -289 3047 -255
rect 3115 -289 3131 -255
rect 3189 -289 3205 -255
rect 3273 -289 3289 -255
rect 3347 -289 3363 -255
rect 3431 -289 3447 -255
rect 3505 -289 3521 -255
rect 3589 -289 3605 -255
rect 3663 -289 3679 -255
rect 3747 -289 3763 -255
rect 3821 -289 3837 -255
rect 3905 -289 3921 -255
rect 3979 -289 3995 -255
rect 4063 -289 4079 -255
rect 4137 -289 4153 -255
rect 4221 -289 4237 -255
rect 4295 -289 4311 -255
rect 4379 -289 4395 -255
rect -4441 -348 -4407 -332
rect -4441 -540 -4407 -524
rect -4283 -348 -4249 -332
rect -4283 -540 -4249 -524
rect -4125 -348 -4091 -332
rect -4125 -540 -4091 -524
rect -3967 -348 -3933 -332
rect -3967 -540 -3933 -524
rect -3809 -348 -3775 -332
rect -3809 -540 -3775 -524
rect -3651 -348 -3617 -332
rect -3651 -540 -3617 -524
rect -3493 -348 -3459 -332
rect -3493 -540 -3459 -524
rect -3335 -348 -3301 -332
rect -3335 -540 -3301 -524
rect -3177 -348 -3143 -332
rect -3177 -540 -3143 -524
rect -3019 -348 -2985 -332
rect -3019 -540 -2985 -524
rect -2861 -348 -2827 -332
rect -2861 -540 -2827 -524
rect -2703 -348 -2669 -332
rect -2703 -540 -2669 -524
rect -2545 -348 -2511 -332
rect -2545 -540 -2511 -524
rect -2387 -348 -2353 -332
rect -2387 -540 -2353 -524
rect -2229 -348 -2195 -332
rect -2229 -540 -2195 -524
rect -2071 -348 -2037 -332
rect -2071 -540 -2037 -524
rect -1913 -348 -1879 -332
rect -1913 -540 -1879 -524
rect -1755 -348 -1721 -332
rect -1755 -540 -1721 -524
rect -1597 -348 -1563 -332
rect -1597 -540 -1563 -524
rect -1439 -348 -1405 -332
rect -1439 -540 -1405 -524
rect -1281 -348 -1247 -332
rect -1281 -540 -1247 -524
rect -1123 -348 -1089 -332
rect -1123 -540 -1089 -524
rect -965 -348 -931 -332
rect -965 -540 -931 -524
rect -807 -348 -773 -332
rect -807 -540 -773 -524
rect -649 -348 -615 -332
rect -649 -540 -615 -524
rect -491 -348 -457 -332
rect -491 -540 -457 -524
rect -333 -348 -299 -332
rect -333 -540 -299 -524
rect -175 -348 -141 -332
rect -175 -540 -141 -524
rect -17 -348 17 -332
rect -17 -540 17 -524
rect 141 -348 175 -332
rect 141 -540 175 -524
rect 299 -348 333 -332
rect 299 -540 333 -524
rect 457 -348 491 -332
rect 457 -540 491 -524
rect 615 -348 649 -332
rect 615 -540 649 -524
rect 773 -348 807 -332
rect 773 -540 807 -524
rect 931 -348 965 -332
rect 931 -540 965 -524
rect 1089 -348 1123 -332
rect 1089 -540 1123 -524
rect 1247 -348 1281 -332
rect 1247 -540 1281 -524
rect 1405 -348 1439 -332
rect 1405 -540 1439 -524
rect 1563 -348 1597 -332
rect 1563 -540 1597 -524
rect 1721 -348 1755 -332
rect 1721 -540 1755 -524
rect 1879 -348 1913 -332
rect 1879 -540 1913 -524
rect 2037 -348 2071 -332
rect 2037 -540 2071 -524
rect 2195 -348 2229 -332
rect 2195 -540 2229 -524
rect 2353 -348 2387 -332
rect 2353 -540 2387 -524
rect 2511 -348 2545 -332
rect 2511 -540 2545 -524
rect 2669 -348 2703 -332
rect 2669 -540 2703 -524
rect 2827 -348 2861 -332
rect 2827 -540 2861 -524
rect 2985 -348 3019 -332
rect 2985 -540 3019 -524
rect 3143 -348 3177 -332
rect 3143 -540 3177 -524
rect 3301 -348 3335 -332
rect 3301 -540 3335 -524
rect 3459 -348 3493 -332
rect 3459 -540 3493 -524
rect 3617 -348 3651 -332
rect 3617 -540 3651 -524
rect 3775 -348 3809 -332
rect 3775 -540 3809 -524
rect 3933 -348 3967 -332
rect 3933 -540 3967 -524
rect 4091 -348 4125 -332
rect 4091 -540 4125 -524
rect 4249 -348 4283 -332
rect 4249 -540 4283 -524
rect 4407 -348 4441 -332
rect 4407 -540 4441 -524
rect -4395 -617 -4379 -583
rect -4311 -617 -4295 -583
rect -4237 -617 -4221 -583
rect -4153 -617 -4137 -583
rect -4079 -617 -4063 -583
rect -3995 -617 -3979 -583
rect -3921 -617 -3905 -583
rect -3837 -617 -3821 -583
rect -3763 -617 -3747 -583
rect -3679 -617 -3663 -583
rect -3605 -617 -3589 -583
rect -3521 -617 -3505 -583
rect -3447 -617 -3431 -583
rect -3363 -617 -3347 -583
rect -3289 -617 -3273 -583
rect -3205 -617 -3189 -583
rect -3131 -617 -3115 -583
rect -3047 -617 -3031 -583
rect -2973 -617 -2957 -583
rect -2889 -617 -2873 -583
rect -2815 -617 -2799 -583
rect -2731 -617 -2715 -583
rect -2657 -617 -2641 -583
rect -2573 -617 -2557 -583
rect -2499 -617 -2483 -583
rect -2415 -617 -2399 -583
rect -2341 -617 -2325 -583
rect -2257 -617 -2241 -583
rect -2183 -617 -2167 -583
rect -2099 -617 -2083 -583
rect -2025 -617 -2009 -583
rect -1941 -617 -1925 -583
rect -1867 -617 -1851 -583
rect -1783 -617 -1767 -583
rect -1709 -617 -1693 -583
rect -1625 -617 -1609 -583
rect -1551 -617 -1535 -583
rect -1467 -617 -1451 -583
rect -1393 -617 -1377 -583
rect -1309 -617 -1293 -583
rect -1235 -617 -1219 -583
rect -1151 -617 -1135 -583
rect -1077 -617 -1061 -583
rect -993 -617 -977 -583
rect -919 -617 -903 -583
rect -835 -617 -819 -583
rect -761 -617 -745 -583
rect -677 -617 -661 -583
rect -603 -617 -587 -583
rect -519 -617 -503 -583
rect -445 -617 -429 -583
rect -361 -617 -345 -583
rect -287 -617 -271 -583
rect -203 -617 -187 -583
rect -129 -617 -113 -583
rect -45 -617 -29 -583
rect 29 -617 45 -583
rect 113 -617 129 -583
rect 187 -617 203 -583
rect 271 -617 287 -583
rect 345 -617 361 -583
rect 429 -617 445 -583
rect 503 -617 519 -583
rect 587 -617 603 -583
rect 661 -617 677 -583
rect 745 -617 761 -583
rect 819 -617 835 -583
rect 903 -617 919 -583
rect 977 -617 993 -583
rect 1061 -617 1077 -583
rect 1135 -617 1151 -583
rect 1219 -617 1235 -583
rect 1293 -617 1309 -583
rect 1377 -617 1393 -583
rect 1451 -617 1467 -583
rect 1535 -617 1551 -583
rect 1609 -617 1625 -583
rect 1693 -617 1709 -583
rect 1767 -617 1783 -583
rect 1851 -617 1867 -583
rect 1925 -617 1941 -583
rect 2009 -617 2025 -583
rect 2083 -617 2099 -583
rect 2167 -617 2183 -583
rect 2241 -617 2257 -583
rect 2325 -617 2341 -583
rect 2399 -617 2415 -583
rect 2483 -617 2499 -583
rect 2557 -617 2573 -583
rect 2641 -617 2657 -583
rect 2715 -617 2731 -583
rect 2799 -617 2815 -583
rect 2873 -617 2889 -583
rect 2957 -617 2973 -583
rect 3031 -617 3047 -583
rect 3115 -617 3131 -583
rect 3189 -617 3205 -583
rect 3273 -617 3289 -583
rect 3347 -617 3363 -583
rect 3431 -617 3447 -583
rect 3505 -617 3521 -583
rect 3589 -617 3605 -583
rect 3663 -617 3679 -583
rect 3747 -617 3763 -583
rect 3821 -617 3837 -583
rect 3905 -617 3921 -583
rect 3979 -617 3995 -583
rect 4063 -617 4079 -583
rect 4137 -617 4153 -583
rect 4221 -617 4237 -583
rect 4295 -617 4311 -583
rect 4379 -617 4395 -583
rect -4395 -725 -4379 -691
rect -4311 -725 -4295 -691
rect -4237 -725 -4221 -691
rect -4153 -725 -4137 -691
rect -4079 -725 -4063 -691
rect -3995 -725 -3979 -691
rect -3921 -725 -3905 -691
rect -3837 -725 -3821 -691
rect -3763 -725 -3747 -691
rect -3679 -725 -3663 -691
rect -3605 -725 -3589 -691
rect -3521 -725 -3505 -691
rect -3447 -725 -3431 -691
rect -3363 -725 -3347 -691
rect -3289 -725 -3273 -691
rect -3205 -725 -3189 -691
rect -3131 -725 -3115 -691
rect -3047 -725 -3031 -691
rect -2973 -725 -2957 -691
rect -2889 -725 -2873 -691
rect -2815 -725 -2799 -691
rect -2731 -725 -2715 -691
rect -2657 -725 -2641 -691
rect -2573 -725 -2557 -691
rect -2499 -725 -2483 -691
rect -2415 -725 -2399 -691
rect -2341 -725 -2325 -691
rect -2257 -725 -2241 -691
rect -2183 -725 -2167 -691
rect -2099 -725 -2083 -691
rect -2025 -725 -2009 -691
rect -1941 -725 -1925 -691
rect -1867 -725 -1851 -691
rect -1783 -725 -1767 -691
rect -1709 -725 -1693 -691
rect -1625 -725 -1609 -691
rect -1551 -725 -1535 -691
rect -1467 -725 -1451 -691
rect -1393 -725 -1377 -691
rect -1309 -725 -1293 -691
rect -1235 -725 -1219 -691
rect -1151 -725 -1135 -691
rect -1077 -725 -1061 -691
rect -993 -725 -977 -691
rect -919 -725 -903 -691
rect -835 -725 -819 -691
rect -761 -725 -745 -691
rect -677 -725 -661 -691
rect -603 -725 -587 -691
rect -519 -725 -503 -691
rect -445 -725 -429 -691
rect -361 -725 -345 -691
rect -287 -725 -271 -691
rect -203 -725 -187 -691
rect -129 -725 -113 -691
rect -45 -725 -29 -691
rect 29 -725 45 -691
rect 113 -725 129 -691
rect 187 -725 203 -691
rect 271 -725 287 -691
rect 345 -725 361 -691
rect 429 -725 445 -691
rect 503 -725 519 -691
rect 587 -725 603 -691
rect 661 -725 677 -691
rect 745 -725 761 -691
rect 819 -725 835 -691
rect 903 -725 919 -691
rect 977 -725 993 -691
rect 1061 -725 1077 -691
rect 1135 -725 1151 -691
rect 1219 -725 1235 -691
rect 1293 -725 1309 -691
rect 1377 -725 1393 -691
rect 1451 -725 1467 -691
rect 1535 -725 1551 -691
rect 1609 -725 1625 -691
rect 1693 -725 1709 -691
rect 1767 -725 1783 -691
rect 1851 -725 1867 -691
rect 1925 -725 1941 -691
rect 2009 -725 2025 -691
rect 2083 -725 2099 -691
rect 2167 -725 2183 -691
rect 2241 -725 2257 -691
rect 2325 -725 2341 -691
rect 2399 -725 2415 -691
rect 2483 -725 2499 -691
rect 2557 -725 2573 -691
rect 2641 -725 2657 -691
rect 2715 -725 2731 -691
rect 2799 -725 2815 -691
rect 2873 -725 2889 -691
rect 2957 -725 2973 -691
rect 3031 -725 3047 -691
rect 3115 -725 3131 -691
rect 3189 -725 3205 -691
rect 3273 -725 3289 -691
rect 3347 -725 3363 -691
rect 3431 -725 3447 -691
rect 3505 -725 3521 -691
rect 3589 -725 3605 -691
rect 3663 -725 3679 -691
rect 3747 -725 3763 -691
rect 3821 -725 3837 -691
rect 3905 -725 3921 -691
rect 3979 -725 3995 -691
rect 4063 -725 4079 -691
rect 4137 -725 4153 -691
rect 4221 -725 4237 -691
rect 4295 -725 4311 -691
rect 4379 -725 4395 -691
rect -4441 -784 -4407 -768
rect -4441 -976 -4407 -960
rect -4283 -784 -4249 -768
rect -4283 -976 -4249 -960
rect -4125 -784 -4091 -768
rect -4125 -976 -4091 -960
rect -3967 -784 -3933 -768
rect -3967 -976 -3933 -960
rect -3809 -784 -3775 -768
rect -3809 -976 -3775 -960
rect -3651 -784 -3617 -768
rect -3651 -976 -3617 -960
rect -3493 -784 -3459 -768
rect -3493 -976 -3459 -960
rect -3335 -784 -3301 -768
rect -3335 -976 -3301 -960
rect -3177 -784 -3143 -768
rect -3177 -976 -3143 -960
rect -3019 -784 -2985 -768
rect -3019 -976 -2985 -960
rect -2861 -784 -2827 -768
rect -2861 -976 -2827 -960
rect -2703 -784 -2669 -768
rect -2703 -976 -2669 -960
rect -2545 -784 -2511 -768
rect -2545 -976 -2511 -960
rect -2387 -784 -2353 -768
rect -2387 -976 -2353 -960
rect -2229 -784 -2195 -768
rect -2229 -976 -2195 -960
rect -2071 -784 -2037 -768
rect -2071 -976 -2037 -960
rect -1913 -784 -1879 -768
rect -1913 -976 -1879 -960
rect -1755 -784 -1721 -768
rect -1755 -976 -1721 -960
rect -1597 -784 -1563 -768
rect -1597 -976 -1563 -960
rect -1439 -784 -1405 -768
rect -1439 -976 -1405 -960
rect -1281 -784 -1247 -768
rect -1281 -976 -1247 -960
rect -1123 -784 -1089 -768
rect -1123 -976 -1089 -960
rect -965 -784 -931 -768
rect -965 -976 -931 -960
rect -807 -784 -773 -768
rect -807 -976 -773 -960
rect -649 -784 -615 -768
rect -649 -976 -615 -960
rect -491 -784 -457 -768
rect -491 -976 -457 -960
rect -333 -784 -299 -768
rect -333 -976 -299 -960
rect -175 -784 -141 -768
rect -175 -976 -141 -960
rect -17 -784 17 -768
rect -17 -976 17 -960
rect 141 -784 175 -768
rect 141 -976 175 -960
rect 299 -784 333 -768
rect 299 -976 333 -960
rect 457 -784 491 -768
rect 457 -976 491 -960
rect 615 -784 649 -768
rect 615 -976 649 -960
rect 773 -784 807 -768
rect 773 -976 807 -960
rect 931 -784 965 -768
rect 931 -976 965 -960
rect 1089 -784 1123 -768
rect 1089 -976 1123 -960
rect 1247 -784 1281 -768
rect 1247 -976 1281 -960
rect 1405 -784 1439 -768
rect 1405 -976 1439 -960
rect 1563 -784 1597 -768
rect 1563 -976 1597 -960
rect 1721 -784 1755 -768
rect 1721 -976 1755 -960
rect 1879 -784 1913 -768
rect 1879 -976 1913 -960
rect 2037 -784 2071 -768
rect 2037 -976 2071 -960
rect 2195 -784 2229 -768
rect 2195 -976 2229 -960
rect 2353 -784 2387 -768
rect 2353 -976 2387 -960
rect 2511 -784 2545 -768
rect 2511 -976 2545 -960
rect 2669 -784 2703 -768
rect 2669 -976 2703 -960
rect 2827 -784 2861 -768
rect 2827 -976 2861 -960
rect 2985 -784 3019 -768
rect 2985 -976 3019 -960
rect 3143 -784 3177 -768
rect 3143 -976 3177 -960
rect 3301 -784 3335 -768
rect 3301 -976 3335 -960
rect 3459 -784 3493 -768
rect 3459 -976 3493 -960
rect 3617 -784 3651 -768
rect 3617 -976 3651 -960
rect 3775 -784 3809 -768
rect 3775 -976 3809 -960
rect 3933 -784 3967 -768
rect 3933 -976 3967 -960
rect 4091 -784 4125 -768
rect 4091 -976 4125 -960
rect 4249 -784 4283 -768
rect 4249 -976 4283 -960
rect 4407 -784 4441 -768
rect 4407 -976 4441 -960
rect -4395 -1053 -4379 -1019
rect -4311 -1053 -4295 -1019
rect -4237 -1053 -4221 -1019
rect -4153 -1053 -4137 -1019
rect -4079 -1053 -4063 -1019
rect -3995 -1053 -3979 -1019
rect -3921 -1053 -3905 -1019
rect -3837 -1053 -3821 -1019
rect -3763 -1053 -3747 -1019
rect -3679 -1053 -3663 -1019
rect -3605 -1053 -3589 -1019
rect -3521 -1053 -3505 -1019
rect -3447 -1053 -3431 -1019
rect -3363 -1053 -3347 -1019
rect -3289 -1053 -3273 -1019
rect -3205 -1053 -3189 -1019
rect -3131 -1053 -3115 -1019
rect -3047 -1053 -3031 -1019
rect -2973 -1053 -2957 -1019
rect -2889 -1053 -2873 -1019
rect -2815 -1053 -2799 -1019
rect -2731 -1053 -2715 -1019
rect -2657 -1053 -2641 -1019
rect -2573 -1053 -2557 -1019
rect -2499 -1053 -2483 -1019
rect -2415 -1053 -2399 -1019
rect -2341 -1053 -2325 -1019
rect -2257 -1053 -2241 -1019
rect -2183 -1053 -2167 -1019
rect -2099 -1053 -2083 -1019
rect -2025 -1053 -2009 -1019
rect -1941 -1053 -1925 -1019
rect -1867 -1053 -1851 -1019
rect -1783 -1053 -1767 -1019
rect -1709 -1053 -1693 -1019
rect -1625 -1053 -1609 -1019
rect -1551 -1053 -1535 -1019
rect -1467 -1053 -1451 -1019
rect -1393 -1053 -1377 -1019
rect -1309 -1053 -1293 -1019
rect -1235 -1053 -1219 -1019
rect -1151 -1053 -1135 -1019
rect -1077 -1053 -1061 -1019
rect -993 -1053 -977 -1019
rect -919 -1053 -903 -1019
rect -835 -1053 -819 -1019
rect -761 -1053 -745 -1019
rect -677 -1053 -661 -1019
rect -603 -1053 -587 -1019
rect -519 -1053 -503 -1019
rect -445 -1053 -429 -1019
rect -361 -1053 -345 -1019
rect -287 -1053 -271 -1019
rect -203 -1053 -187 -1019
rect -129 -1053 -113 -1019
rect -45 -1053 -29 -1019
rect 29 -1053 45 -1019
rect 113 -1053 129 -1019
rect 187 -1053 203 -1019
rect 271 -1053 287 -1019
rect 345 -1053 361 -1019
rect 429 -1053 445 -1019
rect 503 -1053 519 -1019
rect 587 -1053 603 -1019
rect 661 -1053 677 -1019
rect 745 -1053 761 -1019
rect 819 -1053 835 -1019
rect 903 -1053 919 -1019
rect 977 -1053 993 -1019
rect 1061 -1053 1077 -1019
rect 1135 -1053 1151 -1019
rect 1219 -1053 1235 -1019
rect 1293 -1053 1309 -1019
rect 1377 -1053 1393 -1019
rect 1451 -1053 1467 -1019
rect 1535 -1053 1551 -1019
rect 1609 -1053 1625 -1019
rect 1693 -1053 1709 -1019
rect 1767 -1053 1783 -1019
rect 1851 -1053 1867 -1019
rect 1925 -1053 1941 -1019
rect 2009 -1053 2025 -1019
rect 2083 -1053 2099 -1019
rect 2167 -1053 2183 -1019
rect 2241 -1053 2257 -1019
rect 2325 -1053 2341 -1019
rect 2399 -1053 2415 -1019
rect 2483 -1053 2499 -1019
rect 2557 -1053 2573 -1019
rect 2641 -1053 2657 -1019
rect 2715 -1053 2731 -1019
rect 2799 -1053 2815 -1019
rect 2873 -1053 2889 -1019
rect 2957 -1053 2973 -1019
rect 3031 -1053 3047 -1019
rect 3115 -1053 3131 -1019
rect 3189 -1053 3205 -1019
rect 3273 -1053 3289 -1019
rect 3347 -1053 3363 -1019
rect 3431 -1053 3447 -1019
rect 3505 -1053 3521 -1019
rect 3589 -1053 3605 -1019
rect 3663 -1053 3679 -1019
rect 3747 -1053 3763 -1019
rect 3821 -1053 3837 -1019
rect 3905 -1053 3921 -1019
rect 3979 -1053 3995 -1019
rect 4063 -1053 4079 -1019
rect 4137 -1053 4153 -1019
rect 4221 -1053 4237 -1019
rect 4295 -1053 4311 -1019
rect 4379 -1053 4395 -1019
rect -4575 -1157 -4541 -1095
rect 4541 -1157 4575 -1095
rect -4575 -1191 -4479 -1157
rect 4479 -1191 4575 -1157
<< viali >>
rect -4379 1019 -4311 1053
rect -4221 1019 -4153 1053
rect -4063 1019 -3995 1053
rect -3905 1019 -3837 1053
rect -3747 1019 -3679 1053
rect -3589 1019 -3521 1053
rect -3431 1019 -3363 1053
rect -3273 1019 -3205 1053
rect -3115 1019 -3047 1053
rect -2957 1019 -2889 1053
rect -2799 1019 -2731 1053
rect -2641 1019 -2573 1053
rect -2483 1019 -2415 1053
rect -2325 1019 -2257 1053
rect -2167 1019 -2099 1053
rect -2009 1019 -1941 1053
rect -1851 1019 -1783 1053
rect -1693 1019 -1625 1053
rect -1535 1019 -1467 1053
rect -1377 1019 -1309 1053
rect -1219 1019 -1151 1053
rect -1061 1019 -993 1053
rect -903 1019 -835 1053
rect -745 1019 -677 1053
rect -587 1019 -519 1053
rect -429 1019 -361 1053
rect -271 1019 -203 1053
rect -113 1019 -45 1053
rect 45 1019 113 1053
rect 203 1019 271 1053
rect 361 1019 429 1053
rect 519 1019 587 1053
rect 677 1019 745 1053
rect 835 1019 903 1053
rect 993 1019 1061 1053
rect 1151 1019 1219 1053
rect 1309 1019 1377 1053
rect 1467 1019 1535 1053
rect 1625 1019 1693 1053
rect 1783 1019 1851 1053
rect 1941 1019 2009 1053
rect 2099 1019 2167 1053
rect 2257 1019 2325 1053
rect 2415 1019 2483 1053
rect 2573 1019 2641 1053
rect 2731 1019 2799 1053
rect 2889 1019 2957 1053
rect 3047 1019 3115 1053
rect 3205 1019 3273 1053
rect 3363 1019 3431 1053
rect 3521 1019 3589 1053
rect 3679 1019 3747 1053
rect 3837 1019 3905 1053
rect 3995 1019 4063 1053
rect 4153 1019 4221 1053
rect 4311 1019 4379 1053
rect -4441 784 -4407 960
rect -4283 784 -4249 960
rect -4125 784 -4091 960
rect -3967 784 -3933 960
rect -3809 784 -3775 960
rect -3651 784 -3617 960
rect -3493 784 -3459 960
rect -3335 784 -3301 960
rect -3177 784 -3143 960
rect -3019 784 -2985 960
rect -2861 784 -2827 960
rect -2703 784 -2669 960
rect -2545 784 -2511 960
rect -2387 784 -2353 960
rect -2229 784 -2195 960
rect -2071 784 -2037 960
rect -1913 784 -1879 960
rect -1755 784 -1721 960
rect -1597 784 -1563 960
rect -1439 784 -1405 960
rect -1281 784 -1247 960
rect -1123 784 -1089 960
rect -965 784 -931 960
rect -807 784 -773 960
rect -649 784 -615 960
rect -491 784 -457 960
rect -333 784 -299 960
rect -175 784 -141 960
rect -17 784 17 960
rect 141 784 175 960
rect 299 784 333 960
rect 457 784 491 960
rect 615 784 649 960
rect 773 784 807 960
rect 931 784 965 960
rect 1089 784 1123 960
rect 1247 784 1281 960
rect 1405 784 1439 960
rect 1563 784 1597 960
rect 1721 784 1755 960
rect 1879 784 1913 960
rect 2037 784 2071 960
rect 2195 784 2229 960
rect 2353 784 2387 960
rect 2511 784 2545 960
rect 2669 784 2703 960
rect 2827 784 2861 960
rect 2985 784 3019 960
rect 3143 784 3177 960
rect 3301 784 3335 960
rect 3459 784 3493 960
rect 3617 784 3651 960
rect 3775 784 3809 960
rect 3933 784 3967 960
rect 4091 784 4125 960
rect 4249 784 4283 960
rect 4407 784 4441 960
rect -4379 691 -4311 725
rect -4221 691 -4153 725
rect -4063 691 -3995 725
rect -3905 691 -3837 725
rect -3747 691 -3679 725
rect -3589 691 -3521 725
rect -3431 691 -3363 725
rect -3273 691 -3205 725
rect -3115 691 -3047 725
rect -2957 691 -2889 725
rect -2799 691 -2731 725
rect -2641 691 -2573 725
rect -2483 691 -2415 725
rect -2325 691 -2257 725
rect -2167 691 -2099 725
rect -2009 691 -1941 725
rect -1851 691 -1783 725
rect -1693 691 -1625 725
rect -1535 691 -1467 725
rect -1377 691 -1309 725
rect -1219 691 -1151 725
rect -1061 691 -993 725
rect -903 691 -835 725
rect -745 691 -677 725
rect -587 691 -519 725
rect -429 691 -361 725
rect -271 691 -203 725
rect -113 691 -45 725
rect 45 691 113 725
rect 203 691 271 725
rect 361 691 429 725
rect 519 691 587 725
rect 677 691 745 725
rect 835 691 903 725
rect 993 691 1061 725
rect 1151 691 1219 725
rect 1309 691 1377 725
rect 1467 691 1535 725
rect 1625 691 1693 725
rect 1783 691 1851 725
rect 1941 691 2009 725
rect 2099 691 2167 725
rect 2257 691 2325 725
rect 2415 691 2483 725
rect 2573 691 2641 725
rect 2731 691 2799 725
rect 2889 691 2957 725
rect 3047 691 3115 725
rect 3205 691 3273 725
rect 3363 691 3431 725
rect 3521 691 3589 725
rect 3679 691 3747 725
rect 3837 691 3905 725
rect 3995 691 4063 725
rect 4153 691 4221 725
rect 4311 691 4379 725
rect -4379 583 -4311 617
rect -4221 583 -4153 617
rect -4063 583 -3995 617
rect -3905 583 -3837 617
rect -3747 583 -3679 617
rect -3589 583 -3521 617
rect -3431 583 -3363 617
rect -3273 583 -3205 617
rect -3115 583 -3047 617
rect -2957 583 -2889 617
rect -2799 583 -2731 617
rect -2641 583 -2573 617
rect -2483 583 -2415 617
rect -2325 583 -2257 617
rect -2167 583 -2099 617
rect -2009 583 -1941 617
rect -1851 583 -1783 617
rect -1693 583 -1625 617
rect -1535 583 -1467 617
rect -1377 583 -1309 617
rect -1219 583 -1151 617
rect -1061 583 -993 617
rect -903 583 -835 617
rect -745 583 -677 617
rect -587 583 -519 617
rect -429 583 -361 617
rect -271 583 -203 617
rect -113 583 -45 617
rect 45 583 113 617
rect 203 583 271 617
rect 361 583 429 617
rect 519 583 587 617
rect 677 583 745 617
rect 835 583 903 617
rect 993 583 1061 617
rect 1151 583 1219 617
rect 1309 583 1377 617
rect 1467 583 1535 617
rect 1625 583 1693 617
rect 1783 583 1851 617
rect 1941 583 2009 617
rect 2099 583 2167 617
rect 2257 583 2325 617
rect 2415 583 2483 617
rect 2573 583 2641 617
rect 2731 583 2799 617
rect 2889 583 2957 617
rect 3047 583 3115 617
rect 3205 583 3273 617
rect 3363 583 3431 617
rect 3521 583 3589 617
rect 3679 583 3747 617
rect 3837 583 3905 617
rect 3995 583 4063 617
rect 4153 583 4221 617
rect 4311 583 4379 617
rect -4441 348 -4407 524
rect -4283 348 -4249 524
rect -4125 348 -4091 524
rect -3967 348 -3933 524
rect -3809 348 -3775 524
rect -3651 348 -3617 524
rect -3493 348 -3459 524
rect -3335 348 -3301 524
rect -3177 348 -3143 524
rect -3019 348 -2985 524
rect -2861 348 -2827 524
rect -2703 348 -2669 524
rect -2545 348 -2511 524
rect -2387 348 -2353 524
rect -2229 348 -2195 524
rect -2071 348 -2037 524
rect -1913 348 -1879 524
rect -1755 348 -1721 524
rect -1597 348 -1563 524
rect -1439 348 -1405 524
rect -1281 348 -1247 524
rect -1123 348 -1089 524
rect -965 348 -931 524
rect -807 348 -773 524
rect -649 348 -615 524
rect -491 348 -457 524
rect -333 348 -299 524
rect -175 348 -141 524
rect -17 348 17 524
rect 141 348 175 524
rect 299 348 333 524
rect 457 348 491 524
rect 615 348 649 524
rect 773 348 807 524
rect 931 348 965 524
rect 1089 348 1123 524
rect 1247 348 1281 524
rect 1405 348 1439 524
rect 1563 348 1597 524
rect 1721 348 1755 524
rect 1879 348 1913 524
rect 2037 348 2071 524
rect 2195 348 2229 524
rect 2353 348 2387 524
rect 2511 348 2545 524
rect 2669 348 2703 524
rect 2827 348 2861 524
rect 2985 348 3019 524
rect 3143 348 3177 524
rect 3301 348 3335 524
rect 3459 348 3493 524
rect 3617 348 3651 524
rect 3775 348 3809 524
rect 3933 348 3967 524
rect 4091 348 4125 524
rect 4249 348 4283 524
rect 4407 348 4441 524
rect -4379 255 -4311 289
rect -4221 255 -4153 289
rect -4063 255 -3995 289
rect -3905 255 -3837 289
rect -3747 255 -3679 289
rect -3589 255 -3521 289
rect -3431 255 -3363 289
rect -3273 255 -3205 289
rect -3115 255 -3047 289
rect -2957 255 -2889 289
rect -2799 255 -2731 289
rect -2641 255 -2573 289
rect -2483 255 -2415 289
rect -2325 255 -2257 289
rect -2167 255 -2099 289
rect -2009 255 -1941 289
rect -1851 255 -1783 289
rect -1693 255 -1625 289
rect -1535 255 -1467 289
rect -1377 255 -1309 289
rect -1219 255 -1151 289
rect -1061 255 -993 289
rect -903 255 -835 289
rect -745 255 -677 289
rect -587 255 -519 289
rect -429 255 -361 289
rect -271 255 -203 289
rect -113 255 -45 289
rect 45 255 113 289
rect 203 255 271 289
rect 361 255 429 289
rect 519 255 587 289
rect 677 255 745 289
rect 835 255 903 289
rect 993 255 1061 289
rect 1151 255 1219 289
rect 1309 255 1377 289
rect 1467 255 1535 289
rect 1625 255 1693 289
rect 1783 255 1851 289
rect 1941 255 2009 289
rect 2099 255 2167 289
rect 2257 255 2325 289
rect 2415 255 2483 289
rect 2573 255 2641 289
rect 2731 255 2799 289
rect 2889 255 2957 289
rect 3047 255 3115 289
rect 3205 255 3273 289
rect 3363 255 3431 289
rect 3521 255 3589 289
rect 3679 255 3747 289
rect 3837 255 3905 289
rect 3995 255 4063 289
rect 4153 255 4221 289
rect 4311 255 4379 289
rect -4379 147 -4311 181
rect -4221 147 -4153 181
rect -4063 147 -3995 181
rect -3905 147 -3837 181
rect -3747 147 -3679 181
rect -3589 147 -3521 181
rect -3431 147 -3363 181
rect -3273 147 -3205 181
rect -3115 147 -3047 181
rect -2957 147 -2889 181
rect -2799 147 -2731 181
rect -2641 147 -2573 181
rect -2483 147 -2415 181
rect -2325 147 -2257 181
rect -2167 147 -2099 181
rect -2009 147 -1941 181
rect -1851 147 -1783 181
rect -1693 147 -1625 181
rect -1535 147 -1467 181
rect -1377 147 -1309 181
rect -1219 147 -1151 181
rect -1061 147 -993 181
rect -903 147 -835 181
rect -745 147 -677 181
rect -587 147 -519 181
rect -429 147 -361 181
rect -271 147 -203 181
rect -113 147 -45 181
rect 45 147 113 181
rect 203 147 271 181
rect 361 147 429 181
rect 519 147 587 181
rect 677 147 745 181
rect 835 147 903 181
rect 993 147 1061 181
rect 1151 147 1219 181
rect 1309 147 1377 181
rect 1467 147 1535 181
rect 1625 147 1693 181
rect 1783 147 1851 181
rect 1941 147 2009 181
rect 2099 147 2167 181
rect 2257 147 2325 181
rect 2415 147 2483 181
rect 2573 147 2641 181
rect 2731 147 2799 181
rect 2889 147 2957 181
rect 3047 147 3115 181
rect 3205 147 3273 181
rect 3363 147 3431 181
rect 3521 147 3589 181
rect 3679 147 3747 181
rect 3837 147 3905 181
rect 3995 147 4063 181
rect 4153 147 4221 181
rect 4311 147 4379 181
rect -4441 -88 -4407 88
rect -4283 -88 -4249 88
rect -4125 -88 -4091 88
rect -3967 -88 -3933 88
rect -3809 -88 -3775 88
rect -3651 -88 -3617 88
rect -3493 -88 -3459 88
rect -3335 -88 -3301 88
rect -3177 -88 -3143 88
rect -3019 -88 -2985 88
rect -2861 -88 -2827 88
rect -2703 -88 -2669 88
rect -2545 -88 -2511 88
rect -2387 -88 -2353 88
rect -2229 -88 -2195 88
rect -2071 -88 -2037 88
rect -1913 -88 -1879 88
rect -1755 -88 -1721 88
rect -1597 -88 -1563 88
rect -1439 -88 -1405 88
rect -1281 -88 -1247 88
rect -1123 -88 -1089 88
rect -965 -88 -931 88
rect -807 -88 -773 88
rect -649 -88 -615 88
rect -491 -88 -457 88
rect -333 -88 -299 88
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect 299 -88 333 88
rect 457 -88 491 88
rect 615 -88 649 88
rect 773 -88 807 88
rect 931 -88 965 88
rect 1089 -88 1123 88
rect 1247 -88 1281 88
rect 1405 -88 1439 88
rect 1563 -88 1597 88
rect 1721 -88 1755 88
rect 1879 -88 1913 88
rect 2037 -88 2071 88
rect 2195 -88 2229 88
rect 2353 -88 2387 88
rect 2511 -88 2545 88
rect 2669 -88 2703 88
rect 2827 -88 2861 88
rect 2985 -88 3019 88
rect 3143 -88 3177 88
rect 3301 -88 3335 88
rect 3459 -88 3493 88
rect 3617 -88 3651 88
rect 3775 -88 3809 88
rect 3933 -88 3967 88
rect 4091 -88 4125 88
rect 4249 -88 4283 88
rect 4407 -88 4441 88
rect -4379 -181 -4311 -147
rect -4221 -181 -4153 -147
rect -4063 -181 -3995 -147
rect -3905 -181 -3837 -147
rect -3747 -181 -3679 -147
rect -3589 -181 -3521 -147
rect -3431 -181 -3363 -147
rect -3273 -181 -3205 -147
rect -3115 -181 -3047 -147
rect -2957 -181 -2889 -147
rect -2799 -181 -2731 -147
rect -2641 -181 -2573 -147
rect -2483 -181 -2415 -147
rect -2325 -181 -2257 -147
rect -2167 -181 -2099 -147
rect -2009 -181 -1941 -147
rect -1851 -181 -1783 -147
rect -1693 -181 -1625 -147
rect -1535 -181 -1467 -147
rect -1377 -181 -1309 -147
rect -1219 -181 -1151 -147
rect -1061 -181 -993 -147
rect -903 -181 -835 -147
rect -745 -181 -677 -147
rect -587 -181 -519 -147
rect -429 -181 -361 -147
rect -271 -181 -203 -147
rect -113 -181 -45 -147
rect 45 -181 113 -147
rect 203 -181 271 -147
rect 361 -181 429 -147
rect 519 -181 587 -147
rect 677 -181 745 -147
rect 835 -181 903 -147
rect 993 -181 1061 -147
rect 1151 -181 1219 -147
rect 1309 -181 1377 -147
rect 1467 -181 1535 -147
rect 1625 -181 1693 -147
rect 1783 -181 1851 -147
rect 1941 -181 2009 -147
rect 2099 -181 2167 -147
rect 2257 -181 2325 -147
rect 2415 -181 2483 -147
rect 2573 -181 2641 -147
rect 2731 -181 2799 -147
rect 2889 -181 2957 -147
rect 3047 -181 3115 -147
rect 3205 -181 3273 -147
rect 3363 -181 3431 -147
rect 3521 -181 3589 -147
rect 3679 -181 3747 -147
rect 3837 -181 3905 -147
rect 3995 -181 4063 -147
rect 4153 -181 4221 -147
rect 4311 -181 4379 -147
rect -4379 -289 -4311 -255
rect -4221 -289 -4153 -255
rect -4063 -289 -3995 -255
rect -3905 -289 -3837 -255
rect -3747 -289 -3679 -255
rect -3589 -289 -3521 -255
rect -3431 -289 -3363 -255
rect -3273 -289 -3205 -255
rect -3115 -289 -3047 -255
rect -2957 -289 -2889 -255
rect -2799 -289 -2731 -255
rect -2641 -289 -2573 -255
rect -2483 -289 -2415 -255
rect -2325 -289 -2257 -255
rect -2167 -289 -2099 -255
rect -2009 -289 -1941 -255
rect -1851 -289 -1783 -255
rect -1693 -289 -1625 -255
rect -1535 -289 -1467 -255
rect -1377 -289 -1309 -255
rect -1219 -289 -1151 -255
rect -1061 -289 -993 -255
rect -903 -289 -835 -255
rect -745 -289 -677 -255
rect -587 -289 -519 -255
rect -429 -289 -361 -255
rect -271 -289 -203 -255
rect -113 -289 -45 -255
rect 45 -289 113 -255
rect 203 -289 271 -255
rect 361 -289 429 -255
rect 519 -289 587 -255
rect 677 -289 745 -255
rect 835 -289 903 -255
rect 993 -289 1061 -255
rect 1151 -289 1219 -255
rect 1309 -289 1377 -255
rect 1467 -289 1535 -255
rect 1625 -289 1693 -255
rect 1783 -289 1851 -255
rect 1941 -289 2009 -255
rect 2099 -289 2167 -255
rect 2257 -289 2325 -255
rect 2415 -289 2483 -255
rect 2573 -289 2641 -255
rect 2731 -289 2799 -255
rect 2889 -289 2957 -255
rect 3047 -289 3115 -255
rect 3205 -289 3273 -255
rect 3363 -289 3431 -255
rect 3521 -289 3589 -255
rect 3679 -289 3747 -255
rect 3837 -289 3905 -255
rect 3995 -289 4063 -255
rect 4153 -289 4221 -255
rect 4311 -289 4379 -255
rect -4441 -524 -4407 -348
rect -4283 -524 -4249 -348
rect -4125 -524 -4091 -348
rect -3967 -524 -3933 -348
rect -3809 -524 -3775 -348
rect -3651 -524 -3617 -348
rect -3493 -524 -3459 -348
rect -3335 -524 -3301 -348
rect -3177 -524 -3143 -348
rect -3019 -524 -2985 -348
rect -2861 -524 -2827 -348
rect -2703 -524 -2669 -348
rect -2545 -524 -2511 -348
rect -2387 -524 -2353 -348
rect -2229 -524 -2195 -348
rect -2071 -524 -2037 -348
rect -1913 -524 -1879 -348
rect -1755 -524 -1721 -348
rect -1597 -524 -1563 -348
rect -1439 -524 -1405 -348
rect -1281 -524 -1247 -348
rect -1123 -524 -1089 -348
rect -965 -524 -931 -348
rect -807 -524 -773 -348
rect -649 -524 -615 -348
rect -491 -524 -457 -348
rect -333 -524 -299 -348
rect -175 -524 -141 -348
rect -17 -524 17 -348
rect 141 -524 175 -348
rect 299 -524 333 -348
rect 457 -524 491 -348
rect 615 -524 649 -348
rect 773 -524 807 -348
rect 931 -524 965 -348
rect 1089 -524 1123 -348
rect 1247 -524 1281 -348
rect 1405 -524 1439 -348
rect 1563 -524 1597 -348
rect 1721 -524 1755 -348
rect 1879 -524 1913 -348
rect 2037 -524 2071 -348
rect 2195 -524 2229 -348
rect 2353 -524 2387 -348
rect 2511 -524 2545 -348
rect 2669 -524 2703 -348
rect 2827 -524 2861 -348
rect 2985 -524 3019 -348
rect 3143 -524 3177 -348
rect 3301 -524 3335 -348
rect 3459 -524 3493 -348
rect 3617 -524 3651 -348
rect 3775 -524 3809 -348
rect 3933 -524 3967 -348
rect 4091 -524 4125 -348
rect 4249 -524 4283 -348
rect 4407 -524 4441 -348
rect -4379 -617 -4311 -583
rect -4221 -617 -4153 -583
rect -4063 -617 -3995 -583
rect -3905 -617 -3837 -583
rect -3747 -617 -3679 -583
rect -3589 -617 -3521 -583
rect -3431 -617 -3363 -583
rect -3273 -617 -3205 -583
rect -3115 -617 -3047 -583
rect -2957 -617 -2889 -583
rect -2799 -617 -2731 -583
rect -2641 -617 -2573 -583
rect -2483 -617 -2415 -583
rect -2325 -617 -2257 -583
rect -2167 -617 -2099 -583
rect -2009 -617 -1941 -583
rect -1851 -617 -1783 -583
rect -1693 -617 -1625 -583
rect -1535 -617 -1467 -583
rect -1377 -617 -1309 -583
rect -1219 -617 -1151 -583
rect -1061 -617 -993 -583
rect -903 -617 -835 -583
rect -745 -617 -677 -583
rect -587 -617 -519 -583
rect -429 -617 -361 -583
rect -271 -617 -203 -583
rect -113 -617 -45 -583
rect 45 -617 113 -583
rect 203 -617 271 -583
rect 361 -617 429 -583
rect 519 -617 587 -583
rect 677 -617 745 -583
rect 835 -617 903 -583
rect 993 -617 1061 -583
rect 1151 -617 1219 -583
rect 1309 -617 1377 -583
rect 1467 -617 1535 -583
rect 1625 -617 1693 -583
rect 1783 -617 1851 -583
rect 1941 -617 2009 -583
rect 2099 -617 2167 -583
rect 2257 -617 2325 -583
rect 2415 -617 2483 -583
rect 2573 -617 2641 -583
rect 2731 -617 2799 -583
rect 2889 -617 2957 -583
rect 3047 -617 3115 -583
rect 3205 -617 3273 -583
rect 3363 -617 3431 -583
rect 3521 -617 3589 -583
rect 3679 -617 3747 -583
rect 3837 -617 3905 -583
rect 3995 -617 4063 -583
rect 4153 -617 4221 -583
rect 4311 -617 4379 -583
rect -4379 -725 -4311 -691
rect -4221 -725 -4153 -691
rect -4063 -725 -3995 -691
rect -3905 -725 -3837 -691
rect -3747 -725 -3679 -691
rect -3589 -725 -3521 -691
rect -3431 -725 -3363 -691
rect -3273 -725 -3205 -691
rect -3115 -725 -3047 -691
rect -2957 -725 -2889 -691
rect -2799 -725 -2731 -691
rect -2641 -725 -2573 -691
rect -2483 -725 -2415 -691
rect -2325 -725 -2257 -691
rect -2167 -725 -2099 -691
rect -2009 -725 -1941 -691
rect -1851 -725 -1783 -691
rect -1693 -725 -1625 -691
rect -1535 -725 -1467 -691
rect -1377 -725 -1309 -691
rect -1219 -725 -1151 -691
rect -1061 -725 -993 -691
rect -903 -725 -835 -691
rect -745 -725 -677 -691
rect -587 -725 -519 -691
rect -429 -725 -361 -691
rect -271 -725 -203 -691
rect -113 -725 -45 -691
rect 45 -725 113 -691
rect 203 -725 271 -691
rect 361 -725 429 -691
rect 519 -725 587 -691
rect 677 -725 745 -691
rect 835 -725 903 -691
rect 993 -725 1061 -691
rect 1151 -725 1219 -691
rect 1309 -725 1377 -691
rect 1467 -725 1535 -691
rect 1625 -725 1693 -691
rect 1783 -725 1851 -691
rect 1941 -725 2009 -691
rect 2099 -725 2167 -691
rect 2257 -725 2325 -691
rect 2415 -725 2483 -691
rect 2573 -725 2641 -691
rect 2731 -725 2799 -691
rect 2889 -725 2957 -691
rect 3047 -725 3115 -691
rect 3205 -725 3273 -691
rect 3363 -725 3431 -691
rect 3521 -725 3589 -691
rect 3679 -725 3747 -691
rect 3837 -725 3905 -691
rect 3995 -725 4063 -691
rect 4153 -725 4221 -691
rect 4311 -725 4379 -691
rect -4441 -960 -4407 -784
rect -4283 -960 -4249 -784
rect -4125 -960 -4091 -784
rect -3967 -960 -3933 -784
rect -3809 -960 -3775 -784
rect -3651 -960 -3617 -784
rect -3493 -960 -3459 -784
rect -3335 -960 -3301 -784
rect -3177 -960 -3143 -784
rect -3019 -960 -2985 -784
rect -2861 -960 -2827 -784
rect -2703 -960 -2669 -784
rect -2545 -960 -2511 -784
rect -2387 -960 -2353 -784
rect -2229 -960 -2195 -784
rect -2071 -960 -2037 -784
rect -1913 -960 -1879 -784
rect -1755 -960 -1721 -784
rect -1597 -960 -1563 -784
rect -1439 -960 -1405 -784
rect -1281 -960 -1247 -784
rect -1123 -960 -1089 -784
rect -965 -960 -931 -784
rect -807 -960 -773 -784
rect -649 -960 -615 -784
rect -491 -960 -457 -784
rect -333 -960 -299 -784
rect -175 -960 -141 -784
rect -17 -960 17 -784
rect 141 -960 175 -784
rect 299 -960 333 -784
rect 457 -960 491 -784
rect 615 -960 649 -784
rect 773 -960 807 -784
rect 931 -960 965 -784
rect 1089 -960 1123 -784
rect 1247 -960 1281 -784
rect 1405 -960 1439 -784
rect 1563 -960 1597 -784
rect 1721 -960 1755 -784
rect 1879 -960 1913 -784
rect 2037 -960 2071 -784
rect 2195 -960 2229 -784
rect 2353 -960 2387 -784
rect 2511 -960 2545 -784
rect 2669 -960 2703 -784
rect 2827 -960 2861 -784
rect 2985 -960 3019 -784
rect 3143 -960 3177 -784
rect 3301 -960 3335 -784
rect 3459 -960 3493 -784
rect 3617 -960 3651 -784
rect 3775 -960 3809 -784
rect 3933 -960 3967 -784
rect 4091 -960 4125 -784
rect 4249 -960 4283 -784
rect 4407 -960 4441 -784
rect -4379 -1053 -4311 -1019
rect -4221 -1053 -4153 -1019
rect -4063 -1053 -3995 -1019
rect -3905 -1053 -3837 -1019
rect -3747 -1053 -3679 -1019
rect -3589 -1053 -3521 -1019
rect -3431 -1053 -3363 -1019
rect -3273 -1053 -3205 -1019
rect -3115 -1053 -3047 -1019
rect -2957 -1053 -2889 -1019
rect -2799 -1053 -2731 -1019
rect -2641 -1053 -2573 -1019
rect -2483 -1053 -2415 -1019
rect -2325 -1053 -2257 -1019
rect -2167 -1053 -2099 -1019
rect -2009 -1053 -1941 -1019
rect -1851 -1053 -1783 -1019
rect -1693 -1053 -1625 -1019
rect -1535 -1053 -1467 -1019
rect -1377 -1053 -1309 -1019
rect -1219 -1053 -1151 -1019
rect -1061 -1053 -993 -1019
rect -903 -1053 -835 -1019
rect -745 -1053 -677 -1019
rect -587 -1053 -519 -1019
rect -429 -1053 -361 -1019
rect -271 -1053 -203 -1019
rect -113 -1053 -45 -1019
rect 45 -1053 113 -1019
rect 203 -1053 271 -1019
rect 361 -1053 429 -1019
rect 519 -1053 587 -1019
rect 677 -1053 745 -1019
rect 835 -1053 903 -1019
rect 993 -1053 1061 -1019
rect 1151 -1053 1219 -1019
rect 1309 -1053 1377 -1019
rect 1467 -1053 1535 -1019
rect 1625 -1053 1693 -1019
rect 1783 -1053 1851 -1019
rect 1941 -1053 2009 -1019
rect 2099 -1053 2167 -1019
rect 2257 -1053 2325 -1019
rect 2415 -1053 2483 -1019
rect 2573 -1053 2641 -1019
rect 2731 -1053 2799 -1019
rect 2889 -1053 2957 -1019
rect 3047 -1053 3115 -1019
rect 3205 -1053 3273 -1019
rect 3363 -1053 3431 -1019
rect 3521 -1053 3589 -1019
rect 3679 -1053 3747 -1019
rect 3837 -1053 3905 -1019
rect 3995 -1053 4063 -1019
rect 4153 -1053 4221 -1019
rect 4311 -1053 4379 -1019
<< metal1 >>
rect -4391 1053 -4299 1059
rect -4391 1019 -4379 1053
rect -4311 1019 -4299 1053
rect -4391 1013 -4299 1019
rect -4233 1053 -4141 1059
rect -4233 1019 -4221 1053
rect -4153 1019 -4141 1053
rect -4233 1013 -4141 1019
rect -4075 1053 -3983 1059
rect -4075 1019 -4063 1053
rect -3995 1019 -3983 1053
rect -4075 1013 -3983 1019
rect -3917 1053 -3825 1059
rect -3917 1019 -3905 1053
rect -3837 1019 -3825 1053
rect -3917 1013 -3825 1019
rect -3759 1053 -3667 1059
rect -3759 1019 -3747 1053
rect -3679 1019 -3667 1053
rect -3759 1013 -3667 1019
rect -3601 1053 -3509 1059
rect -3601 1019 -3589 1053
rect -3521 1019 -3509 1053
rect -3601 1013 -3509 1019
rect -3443 1053 -3351 1059
rect -3443 1019 -3431 1053
rect -3363 1019 -3351 1053
rect -3443 1013 -3351 1019
rect -3285 1053 -3193 1059
rect -3285 1019 -3273 1053
rect -3205 1019 -3193 1053
rect -3285 1013 -3193 1019
rect -3127 1053 -3035 1059
rect -3127 1019 -3115 1053
rect -3047 1019 -3035 1053
rect -3127 1013 -3035 1019
rect -2969 1053 -2877 1059
rect -2969 1019 -2957 1053
rect -2889 1019 -2877 1053
rect -2969 1013 -2877 1019
rect -2811 1053 -2719 1059
rect -2811 1019 -2799 1053
rect -2731 1019 -2719 1053
rect -2811 1013 -2719 1019
rect -2653 1053 -2561 1059
rect -2653 1019 -2641 1053
rect -2573 1019 -2561 1053
rect -2653 1013 -2561 1019
rect -2495 1053 -2403 1059
rect -2495 1019 -2483 1053
rect -2415 1019 -2403 1053
rect -2495 1013 -2403 1019
rect -2337 1053 -2245 1059
rect -2337 1019 -2325 1053
rect -2257 1019 -2245 1053
rect -2337 1013 -2245 1019
rect -2179 1053 -2087 1059
rect -2179 1019 -2167 1053
rect -2099 1019 -2087 1053
rect -2179 1013 -2087 1019
rect -2021 1053 -1929 1059
rect -2021 1019 -2009 1053
rect -1941 1019 -1929 1053
rect -2021 1013 -1929 1019
rect -1863 1053 -1771 1059
rect -1863 1019 -1851 1053
rect -1783 1019 -1771 1053
rect -1863 1013 -1771 1019
rect -1705 1053 -1613 1059
rect -1705 1019 -1693 1053
rect -1625 1019 -1613 1053
rect -1705 1013 -1613 1019
rect -1547 1053 -1455 1059
rect -1547 1019 -1535 1053
rect -1467 1019 -1455 1053
rect -1547 1013 -1455 1019
rect -1389 1053 -1297 1059
rect -1389 1019 -1377 1053
rect -1309 1019 -1297 1053
rect -1389 1013 -1297 1019
rect -1231 1053 -1139 1059
rect -1231 1019 -1219 1053
rect -1151 1019 -1139 1053
rect -1231 1013 -1139 1019
rect -1073 1053 -981 1059
rect -1073 1019 -1061 1053
rect -993 1019 -981 1053
rect -1073 1013 -981 1019
rect -915 1053 -823 1059
rect -915 1019 -903 1053
rect -835 1019 -823 1053
rect -915 1013 -823 1019
rect -757 1053 -665 1059
rect -757 1019 -745 1053
rect -677 1019 -665 1053
rect -757 1013 -665 1019
rect -599 1053 -507 1059
rect -599 1019 -587 1053
rect -519 1019 -507 1053
rect -599 1013 -507 1019
rect -441 1053 -349 1059
rect -441 1019 -429 1053
rect -361 1019 -349 1053
rect -441 1013 -349 1019
rect -283 1053 -191 1059
rect -283 1019 -271 1053
rect -203 1019 -191 1053
rect -283 1013 -191 1019
rect -125 1053 -33 1059
rect -125 1019 -113 1053
rect -45 1019 -33 1053
rect -125 1013 -33 1019
rect 33 1053 125 1059
rect 33 1019 45 1053
rect 113 1019 125 1053
rect 33 1013 125 1019
rect 191 1053 283 1059
rect 191 1019 203 1053
rect 271 1019 283 1053
rect 191 1013 283 1019
rect 349 1053 441 1059
rect 349 1019 361 1053
rect 429 1019 441 1053
rect 349 1013 441 1019
rect 507 1053 599 1059
rect 507 1019 519 1053
rect 587 1019 599 1053
rect 507 1013 599 1019
rect 665 1053 757 1059
rect 665 1019 677 1053
rect 745 1019 757 1053
rect 665 1013 757 1019
rect 823 1053 915 1059
rect 823 1019 835 1053
rect 903 1019 915 1053
rect 823 1013 915 1019
rect 981 1053 1073 1059
rect 981 1019 993 1053
rect 1061 1019 1073 1053
rect 981 1013 1073 1019
rect 1139 1053 1231 1059
rect 1139 1019 1151 1053
rect 1219 1019 1231 1053
rect 1139 1013 1231 1019
rect 1297 1053 1389 1059
rect 1297 1019 1309 1053
rect 1377 1019 1389 1053
rect 1297 1013 1389 1019
rect 1455 1053 1547 1059
rect 1455 1019 1467 1053
rect 1535 1019 1547 1053
rect 1455 1013 1547 1019
rect 1613 1053 1705 1059
rect 1613 1019 1625 1053
rect 1693 1019 1705 1053
rect 1613 1013 1705 1019
rect 1771 1053 1863 1059
rect 1771 1019 1783 1053
rect 1851 1019 1863 1053
rect 1771 1013 1863 1019
rect 1929 1053 2021 1059
rect 1929 1019 1941 1053
rect 2009 1019 2021 1053
rect 1929 1013 2021 1019
rect 2087 1053 2179 1059
rect 2087 1019 2099 1053
rect 2167 1019 2179 1053
rect 2087 1013 2179 1019
rect 2245 1053 2337 1059
rect 2245 1019 2257 1053
rect 2325 1019 2337 1053
rect 2245 1013 2337 1019
rect 2403 1053 2495 1059
rect 2403 1019 2415 1053
rect 2483 1019 2495 1053
rect 2403 1013 2495 1019
rect 2561 1053 2653 1059
rect 2561 1019 2573 1053
rect 2641 1019 2653 1053
rect 2561 1013 2653 1019
rect 2719 1053 2811 1059
rect 2719 1019 2731 1053
rect 2799 1019 2811 1053
rect 2719 1013 2811 1019
rect 2877 1053 2969 1059
rect 2877 1019 2889 1053
rect 2957 1019 2969 1053
rect 2877 1013 2969 1019
rect 3035 1053 3127 1059
rect 3035 1019 3047 1053
rect 3115 1019 3127 1053
rect 3035 1013 3127 1019
rect 3193 1053 3285 1059
rect 3193 1019 3205 1053
rect 3273 1019 3285 1053
rect 3193 1013 3285 1019
rect 3351 1053 3443 1059
rect 3351 1019 3363 1053
rect 3431 1019 3443 1053
rect 3351 1013 3443 1019
rect 3509 1053 3601 1059
rect 3509 1019 3521 1053
rect 3589 1019 3601 1053
rect 3509 1013 3601 1019
rect 3667 1053 3759 1059
rect 3667 1019 3679 1053
rect 3747 1019 3759 1053
rect 3667 1013 3759 1019
rect 3825 1053 3917 1059
rect 3825 1019 3837 1053
rect 3905 1019 3917 1053
rect 3825 1013 3917 1019
rect 3983 1053 4075 1059
rect 3983 1019 3995 1053
rect 4063 1019 4075 1053
rect 3983 1013 4075 1019
rect 4141 1053 4233 1059
rect 4141 1019 4153 1053
rect 4221 1019 4233 1053
rect 4141 1013 4233 1019
rect 4299 1053 4391 1059
rect 4299 1019 4311 1053
rect 4379 1019 4391 1053
rect 4299 1013 4391 1019
rect -4447 960 -4401 972
rect -4447 784 -4441 960
rect -4407 784 -4401 960
rect -4447 772 -4401 784
rect -4289 960 -4243 972
rect -4289 784 -4283 960
rect -4249 784 -4243 960
rect -4289 772 -4243 784
rect -4131 960 -4085 972
rect -4131 784 -4125 960
rect -4091 784 -4085 960
rect -4131 772 -4085 784
rect -3973 960 -3927 972
rect -3973 784 -3967 960
rect -3933 784 -3927 960
rect -3973 772 -3927 784
rect -3815 960 -3769 972
rect -3815 784 -3809 960
rect -3775 784 -3769 960
rect -3815 772 -3769 784
rect -3657 960 -3611 972
rect -3657 784 -3651 960
rect -3617 784 -3611 960
rect -3657 772 -3611 784
rect -3499 960 -3453 972
rect -3499 784 -3493 960
rect -3459 784 -3453 960
rect -3499 772 -3453 784
rect -3341 960 -3295 972
rect -3341 784 -3335 960
rect -3301 784 -3295 960
rect -3341 772 -3295 784
rect -3183 960 -3137 972
rect -3183 784 -3177 960
rect -3143 784 -3137 960
rect -3183 772 -3137 784
rect -3025 960 -2979 972
rect -3025 784 -3019 960
rect -2985 784 -2979 960
rect -3025 772 -2979 784
rect -2867 960 -2821 972
rect -2867 784 -2861 960
rect -2827 784 -2821 960
rect -2867 772 -2821 784
rect -2709 960 -2663 972
rect -2709 784 -2703 960
rect -2669 784 -2663 960
rect -2709 772 -2663 784
rect -2551 960 -2505 972
rect -2551 784 -2545 960
rect -2511 784 -2505 960
rect -2551 772 -2505 784
rect -2393 960 -2347 972
rect -2393 784 -2387 960
rect -2353 784 -2347 960
rect -2393 772 -2347 784
rect -2235 960 -2189 972
rect -2235 784 -2229 960
rect -2195 784 -2189 960
rect -2235 772 -2189 784
rect -2077 960 -2031 972
rect -2077 784 -2071 960
rect -2037 784 -2031 960
rect -2077 772 -2031 784
rect -1919 960 -1873 972
rect -1919 784 -1913 960
rect -1879 784 -1873 960
rect -1919 772 -1873 784
rect -1761 960 -1715 972
rect -1761 784 -1755 960
rect -1721 784 -1715 960
rect -1761 772 -1715 784
rect -1603 960 -1557 972
rect -1603 784 -1597 960
rect -1563 784 -1557 960
rect -1603 772 -1557 784
rect -1445 960 -1399 972
rect -1445 784 -1439 960
rect -1405 784 -1399 960
rect -1445 772 -1399 784
rect -1287 960 -1241 972
rect -1287 784 -1281 960
rect -1247 784 -1241 960
rect -1287 772 -1241 784
rect -1129 960 -1083 972
rect -1129 784 -1123 960
rect -1089 784 -1083 960
rect -1129 772 -1083 784
rect -971 960 -925 972
rect -971 784 -965 960
rect -931 784 -925 960
rect -971 772 -925 784
rect -813 960 -767 972
rect -813 784 -807 960
rect -773 784 -767 960
rect -813 772 -767 784
rect -655 960 -609 972
rect -655 784 -649 960
rect -615 784 -609 960
rect -655 772 -609 784
rect -497 960 -451 972
rect -497 784 -491 960
rect -457 784 -451 960
rect -497 772 -451 784
rect -339 960 -293 972
rect -339 784 -333 960
rect -299 784 -293 960
rect -339 772 -293 784
rect -181 960 -135 972
rect -181 784 -175 960
rect -141 784 -135 960
rect -181 772 -135 784
rect -23 960 23 972
rect -23 784 -17 960
rect 17 784 23 960
rect -23 772 23 784
rect 135 960 181 972
rect 135 784 141 960
rect 175 784 181 960
rect 135 772 181 784
rect 293 960 339 972
rect 293 784 299 960
rect 333 784 339 960
rect 293 772 339 784
rect 451 960 497 972
rect 451 784 457 960
rect 491 784 497 960
rect 451 772 497 784
rect 609 960 655 972
rect 609 784 615 960
rect 649 784 655 960
rect 609 772 655 784
rect 767 960 813 972
rect 767 784 773 960
rect 807 784 813 960
rect 767 772 813 784
rect 925 960 971 972
rect 925 784 931 960
rect 965 784 971 960
rect 925 772 971 784
rect 1083 960 1129 972
rect 1083 784 1089 960
rect 1123 784 1129 960
rect 1083 772 1129 784
rect 1241 960 1287 972
rect 1241 784 1247 960
rect 1281 784 1287 960
rect 1241 772 1287 784
rect 1399 960 1445 972
rect 1399 784 1405 960
rect 1439 784 1445 960
rect 1399 772 1445 784
rect 1557 960 1603 972
rect 1557 784 1563 960
rect 1597 784 1603 960
rect 1557 772 1603 784
rect 1715 960 1761 972
rect 1715 784 1721 960
rect 1755 784 1761 960
rect 1715 772 1761 784
rect 1873 960 1919 972
rect 1873 784 1879 960
rect 1913 784 1919 960
rect 1873 772 1919 784
rect 2031 960 2077 972
rect 2031 784 2037 960
rect 2071 784 2077 960
rect 2031 772 2077 784
rect 2189 960 2235 972
rect 2189 784 2195 960
rect 2229 784 2235 960
rect 2189 772 2235 784
rect 2347 960 2393 972
rect 2347 784 2353 960
rect 2387 784 2393 960
rect 2347 772 2393 784
rect 2505 960 2551 972
rect 2505 784 2511 960
rect 2545 784 2551 960
rect 2505 772 2551 784
rect 2663 960 2709 972
rect 2663 784 2669 960
rect 2703 784 2709 960
rect 2663 772 2709 784
rect 2821 960 2867 972
rect 2821 784 2827 960
rect 2861 784 2867 960
rect 2821 772 2867 784
rect 2979 960 3025 972
rect 2979 784 2985 960
rect 3019 784 3025 960
rect 2979 772 3025 784
rect 3137 960 3183 972
rect 3137 784 3143 960
rect 3177 784 3183 960
rect 3137 772 3183 784
rect 3295 960 3341 972
rect 3295 784 3301 960
rect 3335 784 3341 960
rect 3295 772 3341 784
rect 3453 960 3499 972
rect 3453 784 3459 960
rect 3493 784 3499 960
rect 3453 772 3499 784
rect 3611 960 3657 972
rect 3611 784 3617 960
rect 3651 784 3657 960
rect 3611 772 3657 784
rect 3769 960 3815 972
rect 3769 784 3775 960
rect 3809 784 3815 960
rect 3769 772 3815 784
rect 3927 960 3973 972
rect 3927 784 3933 960
rect 3967 784 3973 960
rect 3927 772 3973 784
rect 4085 960 4131 972
rect 4085 784 4091 960
rect 4125 784 4131 960
rect 4085 772 4131 784
rect 4243 960 4289 972
rect 4243 784 4249 960
rect 4283 784 4289 960
rect 4243 772 4289 784
rect 4401 960 4447 972
rect 4401 784 4407 960
rect 4441 784 4447 960
rect 4401 772 4447 784
rect -4391 725 -4299 731
rect -4391 691 -4379 725
rect -4311 691 -4299 725
rect -4391 685 -4299 691
rect -4233 725 -4141 731
rect -4233 691 -4221 725
rect -4153 691 -4141 725
rect -4233 685 -4141 691
rect -4075 725 -3983 731
rect -4075 691 -4063 725
rect -3995 691 -3983 725
rect -4075 685 -3983 691
rect -3917 725 -3825 731
rect -3917 691 -3905 725
rect -3837 691 -3825 725
rect -3917 685 -3825 691
rect -3759 725 -3667 731
rect -3759 691 -3747 725
rect -3679 691 -3667 725
rect -3759 685 -3667 691
rect -3601 725 -3509 731
rect -3601 691 -3589 725
rect -3521 691 -3509 725
rect -3601 685 -3509 691
rect -3443 725 -3351 731
rect -3443 691 -3431 725
rect -3363 691 -3351 725
rect -3443 685 -3351 691
rect -3285 725 -3193 731
rect -3285 691 -3273 725
rect -3205 691 -3193 725
rect -3285 685 -3193 691
rect -3127 725 -3035 731
rect -3127 691 -3115 725
rect -3047 691 -3035 725
rect -3127 685 -3035 691
rect -2969 725 -2877 731
rect -2969 691 -2957 725
rect -2889 691 -2877 725
rect -2969 685 -2877 691
rect -2811 725 -2719 731
rect -2811 691 -2799 725
rect -2731 691 -2719 725
rect -2811 685 -2719 691
rect -2653 725 -2561 731
rect -2653 691 -2641 725
rect -2573 691 -2561 725
rect -2653 685 -2561 691
rect -2495 725 -2403 731
rect -2495 691 -2483 725
rect -2415 691 -2403 725
rect -2495 685 -2403 691
rect -2337 725 -2245 731
rect -2337 691 -2325 725
rect -2257 691 -2245 725
rect -2337 685 -2245 691
rect -2179 725 -2087 731
rect -2179 691 -2167 725
rect -2099 691 -2087 725
rect -2179 685 -2087 691
rect -2021 725 -1929 731
rect -2021 691 -2009 725
rect -1941 691 -1929 725
rect -2021 685 -1929 691
rect -1863 725 -1771 731
rect -1863 691 -1851 725
rect -1783 691 -1771 725
rect -1863 685 -1771 691
rect -1705 725 -1613 731
rect -1705 691 -1693 725
rect -1625 691 -1613 725
rect -1705 685 -1613 691
rect -1547 725 -1455 731
rect -1547 691 -1535 725
rect -1467 691 -1455 725
rect -1547 685 -1455 691
rect -1389 725 -1297 731
rect -1389 691 -1377 725
rect -1309 691 -1297 725
rect -1389 685 -1297 691
rect -1231 725 -1139 731
rect -1231 691 -1219 725
rect -1151 691 -1139 725
rect -1231 685 -1139 691
rect -1073 725 -981 731
rect -1073 691 -1061 725
rect -993 691 -981 725
rect -1073 685 -981 691
rect -915 725 -823 731
rect -915 691 -903 725
rect -835 691 -823 725
rect -915 685 -823 691
rect -757 725 -665 731
rect -757 691 -745 725
rect -677 691 -665 725
rect -757 685 -665 691
rect -599 725 -507 731
rect -599 691 -587 725
rect -519 691 -507 725
rect -599 685 -507 691
rect -441 725 -349 731
rect -441 691 -429 725
rect -361 691 -349 725
rect -441 685 -349 691
rect -283 725 -191 731
rect -283 691 -271 725
rect -203 691 -191 725
rect -283 685 -191 691
rect -125 725 -33 731
rect -125 691 -113 725
rect -45 691 -33 725
rect -125 685 -33 691
rect 33 725 125 731
rect 33 691 45 725
rect 113 691 125 725
rect 33 685 125 691
rect 191 725 283 731
rect 191 691 203 725
rect 271 691 283 725
rect 191 685 283 691
rect 349 725 441 731
rect 349 691 361 725
rect 429 691 441 725
rect 349 685 441 691
rect 507 725 599 731
rect 507 691 519 725
rect 587 691 599 725
rect 507 685 599 691
rect 665 725 757 731
rect 665 691 677 725
rect 745 691 757 725
rect 665 685 757 691
rect 823 725 915 731
rect 823 691 835 725
rect 903 691 915 725
rect 823 685 915 691
rect 981 725 1073 731
rect 981 691 993 725
rect 1061 691 1073 725
rect 981 685 1073 691
rect 1139 725 1231 731
rect 1139 691 1151 725
rect 1219 691 1231 725
rect 1139 685 1231 691
rect 1297 725 1389 731
rect 1297 691 1309 725
rect 1377 691 1389 725
rect 1297 685 1389 691
rect 1455 725 1547 731
rect 1455 691 1467 725
rect 1535 691 1547 725
rect 1455 685 1547 691
rect 1613 725 1705 731
rect 1613 691 1625 725
rect 1693 691 1705 725
rect 1613 685 1705 691
rect 1771 725 1863 731
rect 1771 691 1783 725
rect 1851 691 1863 725
rect 1771 685 1863 691
rect 1929 725 2021 731
rect 1929 691 1941 725
rect 2009 691 2021 725
rect 1929 685 2021 691
rect 2087 725 2179 731
rect 2087 691 2099 725
rect 2167 691 2179 725
rect 2087 685 2179 691
rect 2245 725 2337 731
rect 2245 691 2257 725
rect 2325 691 2337 725
rect 2245 685 2337 691
rect 2403 725 2495 731
rect 2403 691 2415 725
rect 2483 691 2495 725
rect 2403 685 2495 691
rect 2561 725 2653 731
rect 2561 691 2573 725
rect 2641 691 2653 725
rect 2561 685 2653 691
rect 2719 725 2811 731
rect 2719 691 2731 725
rect 2799 691 2811 725
rect 2719 685 2811 691
rect 2877 725 2969 731
rect 2877 691 2889 725
rect 2957 691 2969 725
rect 2877 685 2969 691
rect 3035 725 3127 731
rect 3035 691 3047 725
rect 3115 691 3127 725
rect 3035 685 3127 691
rect 3193 725 3285 731
rect 3193 691 3205 725
rect 3273 691 3285 725
rect 3193 685 3285 691
rect 3351 725 3443 731
rect 3351 691 3363 725
rect 3431 691 3443 725
rect 3351 685 3443 691
rect 3509 725 3601 731
rect 3509 691 3521 725
rect 3589 691 3601 725
rect 3509 685 3601 691
rect 3667 725 3759 731
rect 3667 691 3679 725
rect 3747 691 3759 725
rect 3667 685 3759 691
rect 3825 725 3917 731
rect 3825 691 3837 725
rect 3905 691 3917 725
rect 3825 685 3917 691
rect 3983 725 4075 731
rect 3983 691 3995 725
rect 4063 691 4075 725
rect 3983 685 4075 691
rect 4141 725 4233 731
rect 4141 691 4153 725
rect 4221 691 4233 725
rect 4141 685 4233 691
rect 4299 725 4391 731
rect 4299 691 4311 725
rect 4379 691 4391 725
rect 4299 685 4391 691
rect -4391 617 -4299 623
rect -4391 583 -4379 617
rect -4311 583 -4299 617
rect -4391 577 -4299 583
rect -4233 617 -4141 623
rect -4233 583 -4221 617
rect -4153 583 -4141 617
rect -4233 577 -4141 583
rect -4075 617 -3983 623
rect -4075 583 -4063 617
rect -3995 583 -3983 617
rect -4075 577 -3983 583
rect -3917 617 -3825 623
rect -3917 583 -3905 617
rect -3837 583 -3825 617
rect -3917 577 -3825 583
rect -3759 617 -3667 623
rect -3759 583 -3747 617
rect -3679 583 -3667 617
rect -3759 577 -3667 583
rect -3601 617 -3509 623
rect -3601 583 -3589 617
rect -3521 583 -3509 617
rect -3601 577 -3509 583
rect -3443 617 -3351 623
rect -3443 583 -3431 617
rect -3363 583 -3351 617
rect -3443 577 -3351 583
rect -3285 617 -3193 623
rect -3285 583 -3273 617
rect -3205 583 -3193 617
rect -3285 577 -3193 583
rect -3127 617 -3035 623
rect -3127 583 -3115 617
rect -3047 583 -3035 617
rect -3127 577 -3035 583
rect -2969 617 -2877 623
rect -2969 583 -2957 617
rect -2889 583 -2877 617
rect -2969 577 -2877 583
rect -2811 617 -2719 623
rect -2811 583 -2799 617
rect -2731 583 -2719 617
rect -2811 577 -2719 583
rect -2653 617 -2561 623
rect -2653 583 -2641 617
rect -2573 583 -2561 617
rect -2653 577 -2561 583
rect -2495 617 -2403 623
rect -2495 583 -2483 617
rect -2415 583 -2403 617
rect -2495 577 -2403 583
rect -2337 617 -2245 623
rect -2337 583 -2325 617
rect -2257 583 -2245 617
rect -2337 577 -2245 583
rect -2179 617 -2087 623
rect -2179 583 -2167 617
rect -2099 583 -2087 617
rect -2179 577 -2087 583
rect -2021 617 -1929 623
rect -2021 583 -2009 617
rect -1941 583 -1929 617
rect -2021 577 -1929 583
rect -1863 617 -1771 623
rect -1863 583 -1851 617
rect -1783 583 -1771 617
rect -1863 577 -1771 583
rect -1705 617 -1613 623
rect -1705 583 -1693 617
rect -1625 583 -1613 617
rect -1705 577 -1613 583
rect -1547 617 -1455 623
rect -1547 583 -1535 617
rect -1467 583 -1455 617
rect -1547 577 -1455 583
rect -1389 617 -1297 623
rect -1389 583 -1377 617
rect -1309 583 -1297 617
rect -1389 577 -1297 583
rect -1231 617 -1139 623
rect -1231 583 -1219 617
rect -1151 583 -1139 617
rect -1231 577 -1139 583
rect -1073 617 -981 623
rect -1073 583 -1061 617
rect -993 583 -981 617
rect -1073 577 -981 583
rect -915 617 -823 623
rect -915 583 -903 617
rect -835 583 -823 617
rect -915 577 -823 583
rect -757 617 -665 623
rect -757 583 -745 617
rect -677 583 -665 617
rect -757 577 -665 583
rect -599 617 -507 623
rect -599 583 -587 617
rect -519 583 -507 617
rect -599 577 -507 583
rect -441 617 -349 623
rect -441 583 -429 617
rect -361 583 -349 617
rect -441 577 -349 583
rect -283 617 -191 623
rect -283 583 -271 617
rect -203 583 -191 617
rect -283 577 -191 583
rect -125 617 -33 623
rect -125 583 -113 617
rect -45 583 -33 617
rect -125 577 -33 583
rect 33 617 125 623
rect 33 583 45 617
rect 113 583 125 617
rect 33 577 125 583
rect 191 617 283 623
rect 191 583 203 617
rect 271 583 283 617
rect 191 577 283 583
rect 349 617 441 623
rect 349 583 361 617
rect 429 583 441 617
rect 349 577 441 583
rect 507 617 599 623
rect 507 583 519 617
rect 587 583 599 617
rect 507 577 599 583
rect 665 617 757 623
rect 665 583 677 617
rect 745 583 757 617
rect 665 577 757 583
rect 823 617 915 623
rect 823 583 835 617
rect 903 583 915 617
rect 823 577 915 583
rect 981 617 1073 623
rect 981 583 993 617
rect 1061 583 1073 617
rect 981 577 1073 583
rect 1139 617 1231 623
rect 1139 583 1151 617
rect 1219 583 1231 617
rect 1139 577 1231 583
rect 1297 617 1389 623
rect 1297 583 1309 617
rect 1377 583 1389 617
rect 1297 577 1389 583
rect 1455 617 1547 623
rect 1455 583 1467 617
rect 1535 583 1547 617
rect 1455 577 1547 583
rect 1613 617 1705 623
rect 1613 583 1625 617
rect 1693 583 1705 617
rect 1613 577 1705 583
rect 1771 617 1863 623
rect 1771 583 1783 617
rect 1851 583 1863 617
rect 1771 577 1863 583
rect 1929 617 2021 623
rect 1929 583 1941 617
rect 2009 583 2021 617
rect 1929 577 2021 583
rect 2087 617 2179 623
rect 2087 583 2099 617
rect 2167 583 2179 617
rect 2087 577 2179 583
rect 2245 617 2337 623
rect 2245 583 2257 617
rect 2325 583 2337 617
rect 2245 577 2337 583
rect 2403 617 2495 623
rect 2403 583 2415 617
rect 2483 583 2495 617
rect 2403 577 2495 583
rect 2561 617 2653 623
rect 2561 583 2573 617
rect 2641 583 2653 617
rect 2561 577 2653 583
rect 2719 617 2811 623
rect 2719 583 2731 617
rect 2799 583 2811 617
rect 2719 577 2811 583
rect 2877 617 2969 623
rect 2877 583 2889 617
rect 2957 583 2969 617
rect 2877 577 2969 583
rect 3035 617 3127 623
rect 3035 583 3047 617
rect 3115 583 3127 617
rect 3035 577 3127 583
rect 3193 617 3285 623
rect 3193 583 3205 617
rect 3273 583 3285 617
rect 3193 577 3285 583
rect 3351 617 3443 623
rect 3351 583 3363 617
rect 3431 583 3443 617
rect 3351 577 3443 583
rect 3509 617 3601 623
rect 3509 583 3521 617
rect 3589 583 3601 617
rect 3509 577 3601 583
rect 3667 617 3759 623
rect 3667 583 3679 617
rect 3747 583 3759 617
rect 3667 577 3759 583
rect 3825 617 3917 623
rect 3825 583 3837 617
rect 3905 583 3917 617
rect 3825 577 3917 583
rect 3983 617 4075 623
rect 3983 583 3995 617
rect 4063 583 4075 617
rect 3983 577 4075 583
rect 4141 617 4233 623
rect 4141 583 4153 617
rect 4221 583 4233 617
rect 4141 577 4233 583
rect 4299 617 4391 623
rect 4299 583 4311 617
rect 4379 583 4391 617
rect 4299 577 4391 583
rect -4447 524 -4401 536
rect -4447 348 -4441 524
rect -4407 348 -4401 524
rect -4447 336 -4401 348
rect -4289 524 -4243 536
rect -4289 348 -4283 524
rect -4249 348 -4243 524
rect -4289 336 -4243 348
rect -4131 524 -4085 536
rect -4131 348 -4125 524
rect -4091 348 -4085 524
rect -4131 336 -4085 348
rect -3973 524 -3927 536
rect -3973 348 -3967 524
rect -3933 348 -3927 524
rect -3973 336 -3927 348
rect -3815 524 -3769 536
rect -3815 348 -3809 524
rect -3775 348 -3769 524
rect -3815 336 -3769 348
rect -3657 524 -3611 536
rect -3657 348 -3651 524
rect -3617 348 -3611 524
rect -3657 336 -3611 348
rect -3499 524 -3453 536
rect -3499 348 -3493 524
rect -3459 348 -3453 524
rect -3499 336 -3453 348
rect -3341 524 -3295 536
rect -3341 348 -3335 524
rect -3301 348 -3295 524
rect -3341 336 -3295 348
rect -3183 524 -3137 536
rect -3183 348 -3177 524
rect -3143 348 -3137 524
rect -3183 336 -3137 348
rect -3025 524 -2979 536
rect -3025 348 -3019 524
rect -2985 348 -2979 524
rect -3025 336 -2979 348
rect -2867 524 -2821 536
rect -2867 348 -2861 524
rect -2827 348 -2821 524
rect -2867 336 -2821 348
rect -2709 524 -2663 536
rect -2709 348 -2703 524
rect -2669 348 -2663 524
rect -2709 336 -2663 348
rect -2551 524 -2505 536
rect -2551 348 -2545 524
rect -2511 348 -2505 524
rect -2551 336 -2505 348
rect -2393 524 -2347 536
rect -2393 348 -2387 524
rect -2353 348 -2347 524
rect -2393 336 -2347 348
rect -2235 524 -2189 536
rect -2235 348 -2229 524
rect -2195 348 -2189 524
rect -2235 336 -2189 348
rect -2077 524 -2031 536
rect -2077 348 -2071 524
rect -2037 348 -2031 524
rect -2077 336 -2031 348
rect -1919 524 -1873 536
rect -1919 348 -1913 524
rect -1879 348 -1873 524
rect -1919 336 -1873 348
rect -1761 524 -1715 536
rect -1761 348 -1755 524
rect -1721 348 -1715 524
rect -1761 336 -1715 348
rect -1603 524 -1557 536
rect -1603 348 -1597 524
rect -1563 348 -1557 524
rect -1603 336 -1557 348
rect -1445 524 -1399 536
rect -1445 348 -1439 524
rect -1405 348 -1399 524
rect -1445 336 -1399 348
rect -1287 524 -1241 536
rect -1287 348 -1281 524
rect -1247 348 -1241 524
rect -1287 336 -1241 348
rect -1129 524 -1083 536
rect -1129 348 -1123 524
rect -1089 348 -1083 524
rect -1129 336 -1083 348
rect -971 524 -925 536
rect -971 348 -965 524
rect -931 348 -925 524
rect -971 336 -925 348
rect -813 524 -767 536
rect -813 348 -807 524
rect -773 348 -767 524
rect -813 336 -767 348
rect -655 524 -609 536
rect -655 348 -649 524
rect -615 348 -609 524
rect -655 336 -609 348
rect -497 524 -451 536
rect -497 348 -491 524
rect -457 348 -451 524
rect -497 336 -451 348
rect -339 524 -293 536
rect -339 348 -333 524
rect -299 348 -293 524
rect -339 336 -293 348
rect -181 524 -135 536
rect -181 348 -175 524
rect -141 348 -135 524
rect -181 336 -135 348
rect -23 524 23 536
rect -23 348 -17 524
rect 17 348 23 524
rect -23 336 23 348
rect 135 524 181 536
rect 135 348 141 524
rect 175 348 181 524
rect 135 336 181 348
rect 293 524 339 536
rect 293 348 299 524
rect 333 348 339 524
rect 293 336 339 348
rect 451 524 497 536
rect 451 348 457 524
rect 491 348 497 524
rect 451 336 497 348
rect 609 524 655 536
rect 609 348 615 524
rect 649 348 655 524
rect 609 336 655 348
rect 767 524 813 536
rect 767 348 773 524
rect 807 348 813 524
rect 767 336 813 348
rect 925 524 971 536
rect 925 348 931 524
rect 965 348 971 524
rect 925 336 971 348
rect 1083 524 1129 536
rect 1083 348 1089 524
rect 1123 348 1129 524
rect 1083 336 1129 348
rect 1241 524 1287 536
rect 1241 348 1247 524
rect 1281 348 1287 524
rect 1241 336 1287 348
rect 1399 524 1445 536
rect 1399 348 1405 524
rect 1439 348 1445 524
rect 1399 336 1445 348
rect 1557 524 1603 536
rect 1557 348 1563 524
rect 1597 348 1603 524
rect 1557 336 1603 348
rect 1715 524 1761 536
rect 1715 348 1721 524
rect 1755 348 1761 524
rect 1715 336 1761 348
rect 1873 524 1919 536
rect 1873 348 1879 524
rect 1913 348 1919 524
rect 1873 336 1919 348
rect 2031 524 2077 536
rect 2031 348 2037 524
rect 2071 348 2077 524
rect 2031 336 2077 348
rect 2189 524 2235 536
rect 2189 348 2195 524
rect 2229 348 2235 524
rect 2189 336 2235 348
rect 2347 524 2393 536
rect 2347 348 2353 524
rect 2387 348 2393 524
rect 2347 336 2393 348
rect 2505 524 2551 536
rect 2505 348 2511 524
rect 2545 348 2551 524
rect 2505 336 2551 348
rect 2663 524 2709 536
rect 2663 348 2669 524
rect 2703 348 2709 524
rect 2663 336 2709 348
rect 2821 524 2867 536
rect 2821 348 2827 524
rect 2861 348 2867 524
rect 2821 336 2867 348
rect 2979 524 3025 536
rect 2979 348 2985 524
rect 3019 348 3025 524
rect 2979 336 3025 348
rect 3137 524 3183 536
rect 3137 348 3143 524
rect 3177 348 3183 524
rect 3137 336 3183 348
rect 3295 524 3341 536
rect 3295 348 3301 524
rect 3335 348 3341 524
rect 3295 336 3341 348
rect 3453 524 3499 536
rect 3453 348 3459 524
rect 3493 348 3499 524
rect 3453 336 3499 348
rect 3611 524 3657 536
rect 3611 348 3617 524
rect 3651 348 3657 524
rect 3611 336 3657 348
rect 3769 524 3815 536
rect 3769 348 3775 524
rect 3809 348 3815 524
rect 3769 336 3815 348
rect 3927 524 3973 536
rect 3927 348 3933 524
rect 3967 348 3973 524
rect 3927 336 3973 348
rect 4085 524 4131 536
rect 4085 348 4091 524
rect 4125 348 4131 524
rect 4085 336 4131 348
rect 4243 524 4289 536
rect 4243 348 4249 524
rect 4283 348 4289 524
rect 4243 336 4289 348
rect 4401 524 4447 536
rect 4401 348 4407 524
rect 4441 348 4447 524
rect 4401 336 4447 348
rect -4391 289 -4299 295
rect -4391 255 -4379 289
rect -4311 255 -4299 289
rect -4391 249 -4299 255
rect -4233 289 -4141 295
rect -4233 255 -4221 289
rect -4153 255 -4141 289
rect -4233 249 -4141 255
rect -4075 289 -3983 295
rect -4075 255 -4063 289
rect -3995 255 -3983 289
rect -4075 249 -3983 255
rect -3917 289 -3825 295
rect -3917 255 -3905 289
rect -3837 255 -3825 289
rect -3917 249 -3825 255
rect -3759 289 -3667 295
rect -3759 255 -3747 289
rect -3679 255 -3667 289
rect -3759 249 -3667 255
rect -3601 289 -3509 295
rect -3601 255 -3589 289
rect -3521 255 -3509 289
rect -3601 249 -3509 255
rect -3443 289 -3351 295
rect -3443 255 -3431 289
rect -3363 255 -3351 289
rect -3443 249 -3351 255
rect -3285 289 -3193 295
rect -3285 255 -3273 289
rect -3205 255 -3193 289
rect -3285 249 -3193 255
rect -3127 289 -3035 295
rect -3127 255 -3115 289
rect -3047 255 -3035 289
rect -3127 249 -3035 255
rect -2969 289 -2877 295
rect -2969 255 -2957 289
rect -2889 255 -2877 289
rect -2969 249 -2877 255
rect -2811 289 -2719 295
rect -2811 255 -2799 289
rect -2731 255 -2719 289
rect -2811 249 -2719 255
rect -2653 289 -2561 295
rect -2653 255 -2641 289
rect -2573 255 -2561 289
rect -2653 249 -2561 255
rect -2495 289 -2403 295
rect -2495 255 -2483 289
rect -2415 255 -2403 289
rect -2495 249 -2403 255
rect -2337 289 -2245 295
rect -2337 255 -2325 289
rect -2257 255 -2245 289
rect -2337 249 -2245 255
rect -2179 289 -2087 295
rect -2179 255 -2167 289
rect -2099 255 -2087 289
rect -2179 249 -2087 255
rect -2021 289 -1929 295
rect -2021 255 -2009 289
rect -1941 255 -1929 289
rect -2021 249 -1929 255
rect -1863 289 -1771 295
rect -1863 255 -1851 289
rect -1783 255 -1771 289
rect -1863 249 -1771 255
rect -1705 289 -1613 295
rect -1705 255 -1693 289
rect -1625 255 -1613 289
rect -1705 249 -1613 255
rect -1547 289 -1455 295
rect -1547 255 -1535 289
rect -1467 255 -1455 289
rect -1547 249 -1455 255
rect -1389 289 -1297 295
rect -1389 255 -1377 289
rect -1309 255 -1297 289
rect -1389 249 -1297 255
rect -1231 289 -1139 295
rect -1231 255 -1219 289
rect -1151 255 -1139 289
rect -1231 249 -1139 255
rect -1073 289 -981 295
rect -1073 255 -1061 289
rect -993 255 -981 289
rect -1073 249 -981 255
rect -915 289 -823 295
rect -915 255 -903 289
rect -835 255 -823 289
rect -915 249 -823 255
rect -757 289 -665 295
rect -757 255 -745 289
rect -677 255 -665 289
rect -757 249 -665 255
rect -599 289 -507 295
rect -599 255 -587 289
rect -519 255 -507 289
rect -599 249 -507 255
rect -441 289 -349 295
rect -441 255 -429 289
rect -361 255 -349 289
rect -441 249 -349 255
rect -283 289 -191 295
rect -283 255 -271 289
rect -203 255 -191 289
rect -283 249 -191 255
rect -125 289 -33 295
rect -125 255 -113 289
rect -45 255 -33 289
rect -125 249 -33 255
rect 33 289 125 295
rect 33 255 45 289
rect 113 255 125 289
rect 33 249 125 255
rect 191 289 283 295
rect 191 255 203 289
rect 271 255 283 289
rect 191 249 283 255
rect 349 289 441 295
rect 349 255 361 289
rect 429 255 441 289
rect 349 249 441 255
rect 507 289 599 295
rect 507 255 519 289
rect 587 255 599 289
rect 507 249 599 255
rect 665 289 757 295
rect 665 255 677 289
rect 745 255 757 289
rect 665 249 757 255
rect 823 289 915 295
rect 823 255 835 289
rect 903 255 915 289
rect 823 249 915 255
rect 981 289 1073 295
rect 981 255 993 289
rect 1061 255 1073 289
rect 981 249 1073 255
rect 1139 289 1231 295
rect 1139 255 1151 289
rect 1219 255 1231 289
rect 1139 249 1231 255
rect 1297 289 1389 295
rect 1297 255 1309 289
rect 1377 255 1389 289
rect 1297 249 1389 255
rect 1455 289 1547 295
rect 1455 255 1467 289
rect 1535 255 1547 289
rect 1455 249 1547 255
rect 1613 289 1705 295
rect 1613 255 1625 289
rect 1693 255 1705 289
rect 1613 249 1705 255
rect 1771 289 1863 295
rect 1771 255 1783 289
rect 1851 255 1863 289
rect 1771 249 1863 255
rect 1929 289 2021 295
rect 1929 255 1941 289
rect 2009 255 2021 289
rect 1929 249 2021 255
rect 2087 289 2179 295
rect 2087 255 2099 289
rect 2167 255 2179 289
rect 2087 249 2179 255
rect 2245 289 2337 295
rect 2245 255 2257 289
rect 2325 255 2337 289
rect 2245 249 2337 255
rect 2403 289 2495 295
rect 2403 255 2415 289
rect 2483 255 2495 289
rect 2403 249 2495 255
rect 2561 289 2653 295
rect 2561 255 2573 289
rect 2641 255 2653 289
rect 2561 249 2653 255
rect 2719 289 2811 295
rect 2719 255 2731 289
rect 2799 255 2811 289
rect 2719 249 2811 255
rect 2877 289 2969 295
rect 2877 255 2889 289
rect 2957 255 2969 289
rect 2877 249 2969 255
rect 3035 289 3127 295
rect 3035 255 3047 289
rect 3115 255 3127 289
rect 3035 249 3127 255
rect 3193 289 3285 295
rect 3193 255 3205 289
rect 3273 255 3285 289
rect 3193 249 3285 255
rect 3351 289 3443 295
rect 3351 255 3363 289
rect 3431 255 3443 289
rect 3351 249 3443 255
rect 3509 289 3601 295
rect 3509 255 3521 289
rect 3589 255 3601 289
rect 3509 249 3601 255
rect 3667 289 3759 295
rect 3667 255 3679 289
rect 3747 255 3759 289
rect 3667 249 3759 255
rect 3825 289 3917 295
rect 3825 255 3837 289
rect 3905 255 3917 289
rect 3825 249 3917 255
rect 3983 289 4075 295
rect 3983 255 3995 289
rect 4063 255 4075 289
rect 3983 249 4075 255
rect 4141 289 4233 295
rect 4141 255 4153 289
rect 4221 255 4233 289
rect 4141 249 4233 255
rect 4299 289 4391 295
rect 4299 255 4311 289
rect 4379 255 4391 289
rect 4299 249 4391 255
rect -4391 181 -4299 187
rect -4391 147 -4379 181
rect -4311 147 -4299 181
rect -4391 141 -4299 147
rect -4233 181 -4141 187
rect -4233 147 -4221 181
rect -4153 147 -4141 181
rect -4233 141 -4141 147
rect -4075 181 -3983 187
rect -4075 147 -4063 181
rect -3995 147 -3983 181
rect -4075 141 -3983 147
rect -3917 181 -3825 187
rect -3917 147 -3905 181
rect -3837 147 -3825 181
rect -3917 141 -3825 147
rect -3759 181 -3667 187
rect -3759 147 -3747 181
rect -3679 147 -3667 181
rect -3759 141 -3667 147
rect -3601 181 -3509 187
rect -3601 147 -3589 181
rect -3521 147 -3509 181
rect -3601 141 -3509 147
rect -3443 181 -3351 187
rect -3443 147 -3431 181
rect -3363 147 -3351 181
rect -3443 141 -3351 147
rect -3285 181 -3193 187
rect -3285 147 -3273 181
rect -3205 147 -3193 181
rect -3285 141 -3193 147
rect -3127 181 -3035 187
rect -3127 147 -3115 181
rect -3047 147 -3035 181
rect -3127 141 -3035 147
rect -2969 181 -2877 187
rect -2969 147 -2957 181
rect -2889 147 -2877 181
rect -2969 141 -2877 147
rect -2811 181 -2719 187
rect -2811 147 -2799 181
rect -2731 147 -2719 181
rect -2811 141 -2719 147
rect -2653 181 -2561 187
rect -2653 147 -2641 181
rect -2573 147 -2561 181
rect -2653 141 -2561 147
rect -2495 181 -2403 187
rect -2495 147 -2483 181
rect -2415 147 -2403 181
rect -2495 141 -2403 147
rect -2337 181 -2245 187
rect -2337 147 -2325 181
rect -2257 147 -2245 181
rect -2337 141 -2245 147
rect -2179 181 -2087 187
rect -2179 147 -2167 181
rect -2099 147 -2087 181
rect -2179 141 -2087 147
rect -2021 181 -1929 187
rect -2021 147 -2009 181
rect -1941 147 -1929 181
rect -2021 141 -1929 147
rect -1863 181 -1771 187
rect -1863 147 -1851 181
rect -1783 147 -1771 181
rect -1863 141 -1771 147
rect -1705 181 -1613 187
rect -1705 147 -1693 181
rect -1625 147 -1613 181
rect -1705 141 -1613 147
rect -1547 181 -1455 187
rect -1547 147 -1535 181
rect -1467 147 -1455 181
rect -1547 141 -1455 147
rect -1389 181 -1297 187
rect -1389 147 -1377 181
rect -1309 147 -1297 181
rect -1389 141 -1297 147
rect -1231 181 -1139 187
rect -1231 147 -1219 181
rect -1151 147 -1139 181
rect -1231 141 -1139 147
rect -1073 181 -981 187
rect -1073 147 -1061 181
rect -993 147 -981 181
rect -1073 141 -981 147
rect -915 181 -823 187
rect -915 147 -903 181
rect -835 147 -823 181
rect -915 141 -823 147
rect -757 181 -665 187
rect -757 147 -745 181
rect -677 147 -665 181
rect -757 141 -665 147
rect -599 181 -507 187
rect -599 147 -587 181
rect -519 147 -507 181
rect -599 141 -507 147
rect -441 181 -349 187
rect -441 147 -429 181
rect -361 147 -349 181
rect -441 141 -349 147
rect -283 181 -191 187
rect -283 147 -271 181
rect -203 147 -191 181
rect -283 141 -191 147
rect -125 181 -33 187
rect -125 147 -113 181
rect -45 147 -33 181
rect -125 141 -33 147
rect 33 181 125 187
rect 33 147 45 181
rect 113 147 125 181
rect 33 141 125 147
rect 191 181 283 187
rect 191 147 203 181
rect 271 147 283 181
rect 191 141 283 147
rect 349 181 441 187
rect 349 147 361 181
rect 429 147 441 181
rect 349 141 441 147
rect 507 181 599 187
rect 507 147 519 181
rect 587 147 599 181
rect 507 141 599 147
rect 665 181 757 187
rect 665 147 677 181
rect 745 147 757 181
rect 665 141 757 147
rect 823 181 915 187
rect 823 147 835 181
rect 903 147 915 181
rect 823 141 915 147
rect 981 181 1073 187
rect 981 147 993 181
rect 1061 147 1073 181
rect 981 141 1073 147
rect 1139 181 1231 187
rect 1139 147 1151 181
rect 1219 147 1231 181
rect 1139 141 1231 147
rect 1297 181 1389 187
rect 1297 147 1309 181
rect 1377 147 1389 181
rect 1297 141 1389 147
rect 1455 181 1547 187
rect 1455 147 1467 181
rect 1535 147 1547 181
rect 1455 141 1547 147
rect 1613 181 1705 187
rect 1613 147 1625 181
rect 1693 147 1705 181
rect 1613 141 1705 147
rect 1771 181 1863 187
rect 1771 147 1783 181
rect 1851 147 1863 181
rect 1771 141 1863 147
rect 1929 181 2021 187
rect 1929 147 1941 181
rect 2009 147 2021 181
rect 1929 141 2021 147
rect 2087 181 2179 187
rect 2087 147 2099 181
rect 2167 147 2179 181
rect 2087 141 2179 147
rect 2245 181 2337 187
rect 2245 147 2257 181
rect 2325 147 2337 181
rect 2245 141 2337 147
rect 2403 181 2495 187
rect 2403 147 2415 181
rect 2483 147 2495 181
rect 2403 141 2495 147
rect 2561 181 2653 187
rect 2561 147 2573 181
rect 2641 147 2653 181
rect 2561 141 2653 147
rect 2719 181 2811 187
rect 2719 147 2731 181
rect 2799 147 2811 181
rect 2719 141 2811 147
rect 2877 181 2969 187
rect 2877 147 2889 181
rect 2957 147 2969 181
rect 2877 141 2969 147
rect 3035 181 3127 187
rect 3035 147 3047 181
rect 3115 147 3127 181
rect 3035 141 3127 147
rect 3193 181 3285 187
rect 3193 147 3205 181
rect 3273 147 3285 181
rect 3193 141 3285 147
rect 3351 181 3443 187
rect 3351 147 3363 181
rect 3431 147 3443 181
rect 3351 141 3443 147
rect 3509 181 3601 187
rect 3509 147 3521 181
rect 3589 147 3601 181
rect 3509 141 3601 147
rect 3667 181 3759 187
rect 3667 147 3679 181
rect 3747 147 3759 181
rect 3667 141 3759 147
rect 3825 181 3917 187
rect 3825 147 3837 181
rect 3905 147 3917 181
rect 3825 141 3917 147
rect 3983 181 4075 187
rect 3983 147 3995 181
rect 4063 147 4075 181
rect 3983 141 4075 147
rect 4141 181 4233 187
rect 4141 147 4153 181
rect 4221 147 4233 181
rect 4141 141 4233 147
rect 4299 181 4391 187
rect 4299 147 4311 181
rect 4379 147 4391 181
rect 4299 141 4391 147
rect -4447 88 -4401 100
rect -4447 -88 -4441 88
rect -4407 -88 -4401 88
rect -4447 -100 -4401 -88
rect -4289 88 -4243 100
rect -4289 -88 -4283 88
rect -4249 -88 -4243 88
rect -4289 -100 -4243 -88
rect -4131 88 -4085 100
rect -4131 -88 -4125 88
rect -4091 -88 -4085 88
rect -4131 -100 -4085 -88
rect -3973 88 -3927 100
rect -3973 -88 -3967 88
rect -3933 -88 -3927 88
rect -3973 -100 -3927 -88
rect -3815 88 -3769 100
rect -3815 -88 -3809 88
rect -3775 -88 -3769 88
rect -3815 -100 -3769 -88
rect -3657 88 -3611 100
rect -3657 -88 -3651 88
rect -3617 -88 -3611 88
rect -3657 -100 -3611 -88
rect -3499 88 -3453 100
rect -3499 -88 -3493 88
rect -3459 -88 -3453 88
rect -3499 -100 -3453 -88
rect -3341 88 -3295 100
rect -3341 -88 -3335 88
rect -3301 -88 -3295 88
rect -3341 -100 -3295 -88
rect -3183 88 -3137 100
rect -3183 -88 -3177 88
rect -3143 -88 -3137 88
rect -3183 -100 -3137 -88
rect -3025 88 -2979 100
rect -3025 -88 -3019 88
rect -2985 -88 -2979 88
rect -3025 -100 -2979 -88
rect -2867 88 -2821 100
rect -2867 -88 -2861 88
rect -2827 -88 -2821 88
rect -2867 -100 -2821 -88
rect -2709 88 -2663 100
rect -2709 -88 -2703 88
rect -2669 -88 -2663 88
rect -2709 -100 -2663 -88
rect -2551 88 -2505 100
rect -2551 -88 -2545 88
rect -2511 -88 -2505 88
rect -2551 -100 -2505 -88
rect -2393 88 -2347 100
rect -2393 -88 -2387 88
rect -2353 -88 -2347 88
rect -2393 -100 -2347 -88
rect -2235 88 -2189 100
rect -2235 -88 -2229 88
rect -2195 -88 -2189 88
rect -2235 -100 -2189 -88
rect -2077 88 -2031 100
rect -2077 -88 -2071 88
rect -2037 -88 -2031 88
rect -2077 -100 -2031 -88
rect -1919 88 -1873 100
rect -1919 -88 -1913 88
rect -1879 -88 -1873 88
rect -1919 -100 -1873 -88
rect -1761 88 -1715 100
rect -1761 -88 -1755 88
rect -1721 -88 -1715 88
rect -1761 -100 -1715 -88
rect -1603 88 -1557 100
rect -1603 -88 -1597 88
rect -1563 -88 -1557 88
rect -1603 -100 -1557 -88
rect -1445 88 -1399 100
rect -1445 -88 -1439 88
rect -1405 -88 -1399 88
rect -1445 -100 -1399 -88
rect -1287 88 -1241 100
rect -1287 -88 -1281 88
rect -1247 -88 -1241 88
rect -1287 -100 -1241 -88
rect -1129 88 -1083 100
rect -1129 -88 -1123 88
rect -1089 -88 -1083 88
rect -1129 -100 -1083 -88
rect -971 88 -925 100
rect -971 -88 -965 88
rect -931 -88 -925 88
rect -971 -100 -925 -88
rect -813 88 -767 100
rect -813 -88 -807 88
rect -773 -88 -767 88
rect -813 -100 -767 -88
rect -655 88 -609 100
rect -655 -88 -649 88
rect -615 -88 -609 88
rect -655 -100 -609 -88
rect -497 88 -451 100
rect -497 -88 -491 88
rect -457 -88 -451 88
rect -497 -100 -451 -88
rect -339 88 -293 100
rect -339 -88 -333 88
rect -299 -88 -293 88
rect -339 -100 -293 -88
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect 293 88 339 100
rect 293 -88 299 88
rect 333 -88 339 88
rect 293 -100 339 -88
rect 451 88 497 100
rect 451 -88 457 88
rect 491 -88 497 88
rect 451 -100 497 -88
rect 609 88 655 100
rect 609 -88 615 88
rect 649 -88 655 88
rect 609 -100 655 -88
rect 767 88 813 100
rect 767 -88 773 88
rect 807 -88 813 88
rect 767 -100 813 -88
rect 925 88 971 100
rect 925 -88 931 88
rect 965 -88 971 88
rect 925 -100 971 -88
rect 1083 88 1129 100
rect 1083 -88 1089 88
rect 1123 -88 1129 88
rect 1083 -100 1129 -88
rect 1241 88 1287 100
rect 1241 -88 1247 88
rect 1281 -88 1287 88
rect 1241 -100 1287 -88
rect 1399 88 1445 100
rect 1399 -88 1405 88
rect 1439 -88 1445 88
rect 1399 -100 1445 -88
rect 1557 88 1603 100
rect 1557 -88 1563 88
rect 1597 -88 1603 88
rect 1557 -100 1603 -88
rect 1715 88 1761 100
rect 1715 -88 1721 88
rect 1755 -88 1761 88
rect 1715 -100 1761 -88
rect 1873 88 1919 100
rect 1873 -88 1879 88
rect 1913 -88 1919 88
rect 1873 -100 1919 -88
rect 2031 88 2077 100
rect 2031 -88 2037 88
rect 2071 -88 2077 88
rect 2031 -100 2077 -88
rect 2189 88 2235 100
rect 2189 -88 2195 88
rect 2229 -88 2235 88
rect 2189 -100 2235 -88
rect 2347 88 2393 100
rect 2347 -88 2353 88
rect 2387 -88 2393 88
rect 2347 -100 2393 -88
rect 2505 88 2551 100
rect 2505 -88 2511 88
rect 2545 -88 2551 88
rect 2505 -100 2551 -88
rect 2663 88 2709 100
rect 2663 -88 2669 88
rect 2703 -88 2709 88
rect 2663 -100 2709 -88
rect 2821 88 2867 100
rect 2821 -88 2827 88
rect 2861 -88 2867 88
rect 2821 -100 2867 -88
rect 2979 88 3025 100
rect 2979 -88 2985 88
rect 3019 -88 3025 88
rect 2979 -100 3025 -88
rect 3137 88 3183 100
rect 3137 -88 3143 88
rect 3177 -88 3183 88
rect 3137 -100 3183 -88
rect 3295 88 3341 100
rect 3295 -88 3301 88
rect 3335 -88 3341 88
rect 3295 -100 3341 -88
rect 3453 88 3499 100
rect 3453 -88 3459 88
rect 3493 -88 3499 88
rect 3453 -100 3499 -88
rect 3611 88 3657 100
rect 3611 -88 3617 88
rect 3651 -88 3657 88
rect 3611 -100 3657 -88
rect 3769 88 3815 100
rect 3769 -88 3775 88
rect 3809 -88 3815 88
rect 3769 -100 3815 -88
rect 3927 88 3973 100
rect 3927 -88 3933 88
rect 3967 -88 3973 88
rect 3927 -100 3973 -88
rect 4085 88 4131 100
rect 4085 -88 4091 88
rect 4125 -88 4131 88
rect 4085 -100 4131 -88
rect 4243 88 4289 100
rect 4243 -88 4249 88
rect 4283 -88 4289 88
rect 4243 -100 4289 -88
rect 4401 88 4447 100
rect 4401 -88 4407 88
rect 4441 -88 4447 88
rect 4401 -100 4447 -88
rect -4391 -147 -4299 -141
rect -4391 -181 -4379 -147
rect -4311 -181 -4299 -147
rect -4391 -187 -4299 -181
rect -4233 -147 -4141 -141
rect -4233 -181 -4221 -147
rect -4153 -181 -4141 -147
rect -4233 -187 -4141 -181
rect -4075 -147 -3983 -141
rect -4075 -181 -4063 -147
rect -3995 -181 -3983 -147
rect -4075 -187 -3983 -181
rect -3917 -147 -3825 -141
rect -3917 -181 -3905 -147
rect -3837 -181 -3825 -147
rect -3917 -187 -3825 -181
rect -3759 -147 -3667 -141
rect -3759 -181 -3747 -147
rect -3679 -181 -3667 -147
rect -3759 -187 -3667 -181
rect -3601 -147 -3509 -141
rect -3601 -181 -3589 -147
rect -3521 -181 -3509 -147
rect -3601 -187 -3509 -181
rect -3443 -147 -3351 -141
rect -3443 -181 -3431 -147
rect -3363 -181 -3351 -147
rect -3443 -187 -3351 -181
rect -3285 -147 -3193 -141
rect -3285 -181 -3273 -147
rect -3205 -181 -3193 -147
rect -3285 -187 -3193 -181
rect -3127 -147 -3035 -141
rect -3127 -181 -3115 -147
rect -3047 -181 -3035 -147
rect -3127 -187 -3035 -181
rect -2969 -147 -2877 -141
rect -2969 -181 -2957 -147
rect -2889 -181 -2877 -147
rect -2969 -187 -2877 -181
rect -2811 -147 -2719 -141
rect -2811 -181 -2799 -147
rect -2731 -181 -2719 -147
rect -2811 -187 -2719 -181
rect -2653 -147 -2561 -141
rect -2653 -181 -2641 -147
rect -2573 -181 -2561 -147
rect -2653 -187 -2561 -181
rect -2495 -147 -2403 -141
rect -2495 -181 -2483 -147
rect -2415 -181 -2403 -147
rect -2495 -187 -2403 -181
rect -2337 -147 -2245 -141
rect -2337 -181 -2325 -147
rect -2257 -181 -2245 -147
rect -2337 -187 -2245 -181
rect -2179 -147 -2087 -141
rect -2179 -181 -2167 -147
rect -2099 -181 -2087 -147
rect -2179 -187 -2087 -181
rect -2021 -147 -1929 -141
rect -2021 -181 -2009 -147
rect -1941 -181 -1929 -147
rect -2021 -187 -1929 -181
rect -1863 -147 -1771 -141
rect -1863 -181 -1851 -147
rect -1783 -181 -1771 -147
rect -1863 -187 -1771 -181
rect -1705 -147 -1613 -141
rect -1705 -181 -1693 -147
rect -1625 -181 -1613 -147
rect -1705 -187 -1613 -181
rect -1547 -147 -1455 -141
rect -1547 -181 -1535 -147
rect -1467 -181 -1455 -147
rect -1547 -187 -1455 -181
rect -1389 -147 -1297 -141
rect -1389 -181 -1377 -147
rect -1309 -181 -1297 -147
rect -1389 -187 -1297 -181
rect -1231 -147 -1139 -141
rect -1231 -181 -1219 -147
rect -1151 -181 -1139 -147
rect -1231 -187 -1139 -181
rect -1073 -147 -981 -141
rect -1073 -181 -1061 -147
rect -993 -181 -981 -147
rect -1073 -187 -981 -181
rect -915 -147 -823 -141
rect -915 -181 -903 -147
rect -835 -181 -823 -147
rect -915 -187 -823 -181
rect -757 -147 -665 -141
rect -757 -181 -745 -147
rect -677 -181 -665 -147
rect -757 -187 -665 -181
rect -599 -147 -507 -141
rect -599 -181 -587 -147
rect -519 -181 -507 -147
rect -599 -187 -507 -181
rect -441 -147 -349 -141
rect -441 -181 -429 -147
rect -361 -181 -349 -147
rect -441 -187 -349 -181
rect -283 -147 -191 -141
rect -283 -181 -271 -147
rect -203 -181 -191 -147
rect -283 -187 -191 -181
rect -125 -147 -33 -141
rect -125 -181 -113 -147
rect -45 -181 -33 -147
rect -125 -187 -33 -181
rect 33 -147 125 -141
rect 33 -181 45 -147
rect 113 -181 125 -147
rect 33 -187 125 -181
rect 191 -147 283 -141
rect 191 -181 203 -147
rect 271 -181 283 -147
rect 191 -187 283 -181
rect 349 -147 441 -141
rect 349 -181 361 -147
rect 429 -181 441 -147
rect 349 -187 441 -181
rect 507 -147 599 -141
rect 507 -181 519 -147
rect 587 -181 599 -147
rect 507 -187 599 -181
rect 665 -147 757 -141
rect 665 -181 677 -147
rect 745 -181 757 -147
rect 665 -187 757 -181
rect 823 -147 915 -141
rect 823 -181 835 -147
rect 903 -181 915 -147
rect 823 -187 915 -181
rect 981 -147 1073 -141
rect 981 -181 993 -147
rect 1061 -181 1073 -147
rect 981 -187 1073 -181
rect 1139 -147 1231 -141
rect 1139 -181 1151 -147
rect 1219 -181 1231 -147
rect 1139 -187 1231 -181
rect 1297 -147 1389 -141
rect 1297 -181 1309 -147
rect 1377 -181 1389 -147
rect 1297 -187 1389 -181
rect 1455 -147 1547 -141
rect 1455 -181 1467 -147
rect 1535 -181 1547 -147
rect 1455 -187 1547 -181
rect 1613 -147 1705 -141
rect 1613 -181 1625 -147
rect 1693 -181 1705 -147
rect 1613 -187 1705 -181
rect 1771 -147 1863 -141
rect 1771 -181 1783 -147
rect 1851 -181 1863 -147
rect 1771 -187 1863 -181
rect 1929 -147 2021 -141
rect 1929 -181 1941 -147
rect 2009 -181 2021 -147
rect 1929 -187 2021 -181
rect 2087 -147 2179 -141
rect 2087 -181 2099 -147
rect 2167 -181 2179 -147
rect 2087 -187 2179 -181
rect 2245 -147 2337 -141
rect 2245 -181 2257 -147
rect 2325 -181 2337 -147
rect 2245 -187 2337 -181
rect 2403 -147 2495 -141
rect 2403 -181 2415 -147
rect 2483 -181 2495 -147
rect 2403 -187 2495 -181
rect 2561 -147 2653 -141
rect 2561 -181 2573 -147
rect 2641 -181 2653 -147
rect 2561 -187 2653 -181
rect 2719 -147 2811 -141
rect 2719 -181 2731 -147
rect 2799 -181 2811 -147
rect 2719 -187 2811 -181
rect 2877 -147 2969 -141
rect 2877 -181 2889 -147
rect 2957 -181 2969 -147
rect 2877 -187 2969 -181
rect 3035 -147 3127 -141
rect 3035 -181 3047 -147
rect 3115 -181 3127 -147
rect 3035 -187 3127 -181
rect 3193 -147 3285 -141
rect 3193 -181 3205 -147
rect 3273 -181 3285 -147
rect 3193 -187 3285 -181
rect 3351 -147 3443 -141
rect 3351 -181 3363 -147
rect 3431 -181 3443 -147
rect 3351 -187 3443 -181
rect 3509 -147 3601 -141
rect 3509 -181 3521 -147
rect 3589 -181 3601 -147
rect 3509 -187 3601 -181
rect 3667 -147 3759 -141
rect 3667 -181 3679 -147
rect 3747 -181 3759 -147
rect 3667 -187 3759 -181
rect 3825 -147 3917 -141
rect 3825 -181 3837 -147
rect 3905 -181 3917 -147
rect 3825 -187 3917 -181
rect 3983 -147 4075 -141
rect 3983 -181 3995 -147
rect 4063 -181 4075 -147
rect 3983 -187 4075 -181
rect 4141 -147 4233 -141
rect 4141 -181 4153 -147
rect 4221 -181 4233 -147
rect 4141 -187 4233 -181
rect 4299 -147 4391 -141
rect 4299 -181 4311 -147
rect 4379 -181 4391 -147
rect 4299 -187 4391 -181
rect -4391 -255 -4299 -249
rect -4391 -289 -4379 -255
rect -4311 -289 -4299 -255
rect -4391 -295 -4299 -289
rect -4233 -255 -4141 -249
rect -4233 -289 -4221 -255
rect -4153 -289 -4141 -255
rect -4233 -295 -4141 -289
rect -4075 -255 -3983 -249
rect -4075 -289 -4063 -255
rect -3995 -289 -3983 -255
rect -4075 -295 -3983 -289
rect -3917 -255 -3825 -249
rect -3917 -289 -3905 -255
rect -3837 -289 -3825 -255
rect -3917 -295 -3825 -289
rect -3759 -255 -3667 -249
rect -3759 -289 -3747 -255
rect -3679 -289 -3667 -255
rect -3759 -295 -3667 -289
rect -3601 -255 -3509 -249
rect -3601 -289 -3589 -255
rect -3521 -289 -3509 -255
rect -3601 -295 -3509 -289
rect -3443 -255 -3351 -249
rect -3443 -289 -3431 -255
rect -3363 -289 -3351 -255
rect -3443 -295 -3351 -289
rect -3285 -255 -3193 -249
rect -3285 -289 -3273 -255
rect -3205 -289 -3193 -255
rect -3285 -295 -3193 -289
rect -3127 -255 -3035 -249
rect -3127 -289 -3115 -255
rect -3047 -289 -3035 -255
rect -3127 -295 -3035 -289
rect -2969 -255 -2877 -249
rect -2969 -289 -2957 -255
rect -2889 -289 -2877 -255
rect -2969 -295 -2877 -289
rect -2811 -255 -2719 -249
rect -2811 -289 -2799 -255
rect -2731 -289 -2719 -255
rect -2811 -295 -2719 -289
rect -2653 -255 -2561 -249
rect -2653 -289 -2641 -255
rect -2573 -289 -2561 -255
rect -2653 -295 -2561 -289
rect -2495 -255 -2403 -249
rect -2495 -289 -2483 -255
rect -2415 -289 -2403 -255
rect -2495 -295 -2403 -289
rect -2337 -255 -2245 -249
rect -2337 -289 -2325 -255
rect -2257 -289 -2245 -255
rect -2337 -295 -2245 -289
rect -2179 -255 -2087 -249
rect -2179 -289 -2167 -255
rect -2099 -289 -2087 -255
rect -2179 -295 -2087 -289
rect -2021 -255 -1929 -249
rect -2021 -289 -2009 -255
rect -1941 -289 -1929 -255
rect -2021 -295 -1929 -289
rect -1863 -255 -1771 -249
rect -1863 -289 -1851 -255
rect -1783 -289 -1771 -255
rect -1863 -295 -1771 -289
rect -1705 -255 -1613 -249
rect -1705 -289 -1693 -255
rect -1625 -289 -1613 -255
rect -1705 -295 -1613 -289
rect -1547 -255 -1455 -249
rect -1547 -289 -1535 -255
rect -1467 -289 -1455 -255
rect -1547 -295 -1455 -289
rect -1389 -255 -1297 -249
rect -1389 -289 -1377 -255
rect -1309 -289 -1297 -255
rect -1389 -295 -1297 -289
rect -1231 -255 -1139 -249
rect -1231 -289 -1219 -255
rect -1151 -289 -1139 -255
rect -1231 -295 -1139 -289
rect -1073 -255 -981 -249
rect -1073 -289 -1061 -255
rect -993 -289 -981 -255
rect -1073 -295 -981 -289
rect -915 -255 -823 -249
rect -915 -289 -903 -255
rect -835 -289 -823 -255
rect -915 -295 -823 -289
rect -757 -255 -665 -249
rect -757 -289 -745 -255
rect -677 -289 -665 -255
rect -757 -295 -665 -289
rect -599 -255 -507 -249
rect -599 -289 -587 -255
rect -519 -289 -507 -255
rect -599 -295 -507 -289
rect -441 -255 -349 -249
rect -441 -289 -429 -255
rect -361 -289 -349 -255
rect -441 -295 -349 -289
rect -283 -255 -191 -249
rect -283 -289 -271 -255
rect -203 -289 -191 -255
rect -283 -295 -191 -289
rect -125 -255 -33 -249
rect -125 -289 -113 -255
rect -45 -289 -33 -255
rect -125 -295 -33 -289
rect 33 -255 125 -249
rect 33 -289 45 -255
rect 113 -289 125 -255
rect 33 -295 125 -289
rect 191 -255 283 -249
rect 191 -289 203 -255
rect 271 -289 283 -255
rect 191 -295 283 -289
rect 349 -255 441 -249
rect 349 -289 361 -255
rect 429 -289 441 -255
rect 349 -295 441 -289
rect 507 -255 599 -249
rect 507 -289 519 -255
rect 587 -289 599 -255
rect 507 -295 599 -289
rect 665 -255 757 -249
rect 665 -289 677 -255
rect 745 -289 757 -255
rect 665 -295 757 -289
rect 823 -255 915 -249
rect 823 -289 835 -255
rect 903 -289 915 -255
rect 823 -295 915 -289
rect 981 -255 1073 -249
rect 981 -289 993 -255
rect 1061 -289 1073 -255
rect 981 -295 1073 -289
rect 1139 -255 1231 -249
rect 1139 -289 1151 -255
rect 1219 -289 1231 -255
rect 1139 -295 1231 -289
rect 1297 -255 1389 -249
rect 1297 -289 1309 -255
rect 1377 -289 1389 -255
rect 1297 -295 1389 -289
rect 1455 -255 1547 -249
rect 1455 -289 1467 -255
rect 1535 -289 1547 -255
rect 1455 -295 1547 -289
rect 1613 -255 1705 -249
rect 1613 -289 1625 -255
rect 1693 -289 1705 -255
rect 1613 -295 1705 -289
rect 1771 -255 1863 -249
rect 1771 -289 1783 -255
rect 1851 -289 1863 -255
rect 1771 -295 1863 -289
rect 1929 -255 2021 -249
rect 1929 -289 1941 -255
rect 2009 -289 2021 -255
rect 1929 -295 2021 -289
rect 2087 -255 2179 -249
rect 2087 -289 2099 -255
rect 2167 -289 2179 -255
rect 2087 -295 2179 -289
rect 2245 -255 2337 -249
rect 2245 -289 2257 -255
rect 2325 -289 2337 -255
rect 2245 -295 2337 -289
rect 2403 -255 2495 -249
rect 2403 -289 2415 -255
rect 2483 -289 2495 -255
rect 2403 -295 2495 -289
rect 2561 -255 2653 -249
rect 2561 -289 2573 -255
rect 2641 -289 2653 -255
rect 2561 -295 2653 -289
rect 2719 -255 2811 -249
rect 2719 -289 2731 -255
rect 2799 -289 2811 -255
rect 2719 -295 2811 -289
rect 2877 -255 2969 -249
rect 2877 -289 2889 -255
rect 2957 -289 2969 -255
rect 2877 -295 2969 -289
rect 3035 -255 3127 -249
rect 3035 -289 3047 -255
rect 3115 -289 3127 -255
rect 3035 -295 3127 -289
rect 3193 -255 3285 -249
rect 3193 -289 3205 -255
rect 3273 -289 3285 -255
rect 3193 -295 3285 -289
rect 3351 -255 3443 -249
rect 3351 -289 3363 -255
rect 3431 -289 3443 -255
rect 3351 -295 3443 -289
rect 3509 -255 3601 -249
rect 3509 -289 3521 -255
rect 3589 -289 3601 -255
rect 3509 -295 3601 -289
rect 3667 -255 3759 -249
rect 3667 -289 3679 -255
rect 3747 -289 3759 -255
rect 3667 -295 3759 -289
rect 3825 -255 3917 -249
rect 3825 -289 3837 -255
rect 3905 -289 3917 -255
rect 3825 -295 3917 -289
rect 3983 -255 4075 -249
rect 3983 -289 3995 -255
rect 4063 -289 4075 -255
rect 3983 -295 4075 -289
rect 4141 -255 4233 -249
rect 4141 -289 4153 -255
rect 4221 -289 4233 -255
rect 4141 -295 4233 -289
rect 4299 -255 4391 -249
rect 4299 -289 4311 -255
rect 4379 -289 4391 -255
rect 4299 -295 4391 -289
rect -4447 -348 -4401 -336
rect -4447 -524 -4441 -348
rect -4407 -524 -4401 -348
rect -4447 -536 -4401 -524
rect -4289 -348 -4243 -336
rect -4289 -524 -4283 -348
rect -4249 -524 -4243 -348
rect -4289 -536 -4243 -524
rect -4131 -348 -4085 -336
rect -4131 -524 -4125 -348
rect -4091 -524 -4085 -348
rect -4131 -536 -4085 -524
rect -3973 -348 -3927 -336
rect -3973 -524 -3967 -348
rect -3933 -524 -3927 -348
rect -3973 -536 -3927 -524
rect -3815 -348 -3769 -336
rect -3815 -524 -3809 -348
rect -3775 -524 -3769 -348
rect -3815 -536 -3769 -524
rect -3657 -348 -3611 -336
rect -3657 -524 -3651 -348
rect -3617 -524 -3611 -348
rect -3657 -536 -3611 -524
rect -3499 -348 -3453 -336
rect -3499 -524 -3493 -348
rect -3459 -524 -3453 -348
rect -3499 -536 -3453 -524
rect -3341 -348 -3295 -336
rect -3341 -524 -3335 -348
rect -3301 -524 -3295 -348
rect -3341 -536 -3295 -524
rect -3183 -348 -3137 -336
rect -3183 -524 -3177 -348
rect -3143 -524 -3137 -348
rect -3183 -536 -3137 -524
rect -3025 -348 -2979 -336
rect -3025 -524 -3019 -348
rect -2985 -524 -2979 -348
rect -3025 -536 -2979 -524
rect -2867 -348 -2821 -336
rect -2867 -524 -2861 -348
rect -2827 -524 -2821 -348
rect -2867 -536 -2821 -524
rect -2709 -348 -2663 -336
rect -2709 -524 -2703 -348
rect -2669 -524 -2663 -348
rect -2709 -536 -2663 -524
rect -2551 -348 -2505 -336
rect -2551 -524 -2545 -348
rect -2511 -524 -2505 -348
rect -2551 -536 -2505 -524
rect -2393 -348 -2347 -336
rect -2393 -524 -2387 -348
rect -2353 -524 -2347 -348
rect -2393 -536 -2347 -524
rect -2235 -348 -2189 -336
rect -2235 -524 -2229 -348
rect -2195 -524 -2189 -348
rect -2235 -536 -2189 -524
rect -2077 -348 -2031 -336
rect -2077 -524 -2071 -348
rect -2037 -524 -2031 -348
rect -2077 -536 -2031 -524
rect -1919 -348 -1873 -336
rect -1919 -524 -1913 -348
rect -1879 -524 -1873 -348
rect -1919 -536 -1873 -524
rect -1761 -348 -1715 -336
rect -1761 -524 -1755 -348
rect -1721 -524 -1715 -348
rect -1761 -536 -1715 -524
rect -1603 -348 -1557 -336
rect -1603 -524 -1597 -348
rect -1563 -524 -1557 -348
rect -1603 -536 -1557 -524
rect -1445 -348 -1399 -336
rect -1445 -524 -1439 -348
rect -1405 -524 -1399 -348
rect -1445 -536 -1399 -524
rect -1287 -348 -1241 -336
rect -1287 -524 -1281 -348
rect -1247 -524 -1241 -348
rect -1287 -536 -1241 -524
rect -1129 -348 -1083 -336
rect -1129 -524 -1123 -348
rect -1089 -524 -1083 -348
rect -1129 -536 -1083 -524
rect -971 -348 -925 -336
rect -971 -524 -965 -348
rect -931 -524 -925 -348
rect -971 -536 -925 -524
rect -813 -348 -767 -336
rect -813 -524 -807 -348
rect -773 -524 -767 -348
rect -813 -536 -767 -524
rect -655 -348 -609 -336
rect -655 -524 -649 -348
rect -615 -524 -609 -348
rect -655 -536 -609 -524
rect -497 -348 -451 -336
rect -497 -524 -491 -348
rect -457 -524 -451 -348
rect -497 -536 -451 -524
rect -339 -348 -293 -336
rect -339 -524 -333 -348
rect -299 -524 -293 -348
rect -339 -536 -293 -524
rect -181 -348 -135 -336
rect -181 -524 -175 -348
rect -141 -524 -135 -348
rect -181 -536 -135 -524
rect -23 -348 23 -336
rect -23 -524 -17 -348
rect 17 -524 23 -348
rect -23 -536 23 -524
rect 135 -348 181 -336
rect 135 -524 141 -348
rect 175 -524 181 -348
rect 135 -536 181 -524
rect 293 -348 339 -336
rect 293 -524 299 -348
rect 333 -524 339 -348
rect 293 -536 339 -524
rect 451 -348 497 -336
rect 451 -524 457 -348
rect 491 -524 497 -348
rect 451 -536 497 -524
rect 609 -348 655 -336
rect 609 -524 615 -348
rect 649 -524 655 -348
rect 609 -536 655 -524
rect 767 -348 813 -336
rect 767 -524 773 -348
rect 807 -524 813 -348
rect 767 -536 813 -524
rect 925 -348 971 -336
rect 925 -524 931 -348
rect 965 -524 971 -348
rect 925 -536 971 -524
rect 1083 -348 1129 -336
rect 1083 -524 1089 -348
rect 1123 -524 1129 -348
rect 1083 -536 1129 -524
rect 1241 -348 1287 -336
rect 1241 -524 1247 -348
rect 1281 -524 1287 -348
rect 1241 -536 1287 -524
rect 1399 -348 1445 -336
rect 1399 -524 1405 -348
rect 1439 -524 1445 -348
rect 1399 -536 1445 -524
rect 1557 -348 1603 -336
rect 1557 -524 1563 -348
rect 1597 -524 1603 -348
rect 1557 -536 1603 -524
rect 1715 -348 1761 -336
rect 1715 -524 1721 -348
rect 1755 -524 1761 -348
rect 1715 -536 1761 -524
rect 1873 -348 1919 -336
rect 1873 -524 1879 -348
rect 1913 -524 1919 -348
rect 1873 -536 1919 -524
rect 2031 -348 2077 -336
rect 2031 -524 2037 -348
rect 2071 -524 2077 -348
rect 2031 -536 2077 -524
rect 2189 -348 2235 -336
rect 2189 -524 2195 -348
rect 2229 -524 2235 -348
rect 2189 -536 2235 -524
rect 2347 -348 2393 -336
rect 2347 -524 2353 -348
rect 2387 -524 2393 -348
rect 2347 -536 2393 -524
rect 2505 -348 2551 -336
rect 2505 -524 2511 -348
rect 2545 -524 2551 -348
rect 2505 -536 2551 -524
rect 2663 -348 2709 -336
rect 2663 -524 2669 -348
rect 2703 -524 2709 -348
rect 2663 -536 2709 -524
rect 2821 -348 2867 -336
rect 2821 -524 2827 -348
rect 2861 -524 2867 -348
rect 2821 -536 2867 -524
rect 2979 -348 3025 -336
rect 2979 -524 2985 -348
rect 3019 -524 3025 -348
rect 2979 -536 3025 -524
rect 3137 -348 3183 -336
rect 3137 -524 3143 -348
rect 3177 -524 3183 -348
rect 3137 -536 3183 -524
rect 3295 -348 3341 -336
rect 3295 -524 3301 -348
rect 3335 -524 3341 -348
rect 3295 -536 3341 -524
rect 3453 -348 3499 -336
rect 3453 -524 3459 -348
rect 3493 -524 3499 -348
rect 3453 -536 3499 -524
rect 3611 -348 3657 -336
rect 3611 -524 3617 -348
rect 3651 -524 3657 -348
rect 3611 -536 3657 -524
rect 3769 -348 3815 -336
rect 3769 -524 3775 -348
rect 3809 -524 3815 -348
rect 3769 -536 3815 -524
rect 3927 -348 3973 -336
rect 3927 -524 3933 -348
rect 3967 -524 3973 -348
rect 3927 -536 3973 -524
rect 4085 -348 4131 -336
rect 4085 -524 4091 -348
rect 4125 -524 4131 -348
rect 4085 -536 4131 -524
rect 4243 -348 4289 -336
rect 4243 -524 4249 -348
rect 4283 -524 4289 -348
rect 4243 -536 4289 -524
rect 4401 -348 4447 -336
rect 4401 -524 4407 -348
rect 4441 -524 4447 -348
rect 4401 -536 4447 -524
rect -4391 -583 -4299 -577
rect -4391 -617 -4379 -583
rect -4311 -617 -4299 -583
rect -4391 -623 -4299 -617
rect -4233 -583 -4141 -577
rect -4233 -617 -4221 -583
rect -4153 -617 -4141 -583
rect -4233 -623 -4141 -617
rect -4075 -583 -3983 -577
rect -4075 -617 -4063 -583
rect -3995 -617 -3983 -583
rect -4075 -623 -3983 -617
rect -3917 -583 -3825 -577
rect -3917 -617 -3905 -583
rect -3837 -617 -3825 -583
rect -3917 -623 -3825 -617
rect -3759 -583 -3667 -577
rect -3759 -617 -3747 -583
rect -3679 -617 -3667 -583
rect -3759 -623 -3667 -617
rect -3601 -583 -3509 -577
rect -3601 -617 -3589 -583
rect -3521 -617 -3509 -583
rect -3601 -623 -3509 -617
rect -3443 -583 -3351 -577
rect -3443 -617 -3431 -583
rect -3363 -617 -3351 -583
rect -3443 -623 -3351 -617
rect -3285 -583 -3193 -577
rect -3285 -617 -3273 -583
rect -3205 -617 -3193 -583
rect -3285 -623 -3193 -617
rect -3127 -583 -3035 -577
rect -3127 -617 -3115 -583
rect -3047 -617 -3035 -583
rect -3127 -623 -3035 -617
rect -2969 -583 -2877 -577
rect -2969 -617 -2957 -583
rect -2889 -617 -2877 -583
rect -2969 -623 -2877 -617
rect -2811 -583 -2719 -577
rect -2811 -617 -2799 -583
rect -2731 -617 -2719 -583
rect -2811 -623 -2719 -617
rect -2653 -583 -2561 -577
rect -2653 -617 -2641 -583
rect -2573 -617 -2561 -583
rect -2653 -623 -2561 -617
rect -2495 -583 -2403 -577
rect -2495 -617 -2483 -583
rect -2415 -617 -2403 -583
rect -2495 -623 -2403 -617
rect -2337 -583 -2245 -577
rect -2337 -617 -2325 -583
rect -2257 -617 -2245 -583
rect -2337 -623 -2245 -617
rect -2179 -583 -2087 -577
rect -2179 -617 -2167 -583
rect -2099 -617 -2087 -583
rect -2179 -623 -2087 -617
rect -2021 -583 -1929 -577
rect -2021 -617 -2009 -583
rect -1941 -617 -1929 -583
rect -2021 -623 -1929 -617
rect -1863 -583 -1771 -577
rect -1863 -617 -1851 -583
rect -1783 -617 -1771 -583
rect -1863 -623 -1771 -617
rect -1705 -583 -1613 -577
rect -1705 -617 -1693 -583
rect -1625 -617 -1613 -583
rect -1705 -623 -1613 -617
rect -1547 -583 -1455 -577
rect -1547 -617 -1535 -583
rect -1467 -617 -1455 -583
rect -1547 -623 -1455 -617
rect -1389 -583 -1297 -577
rect -1389 -617 -1377 -583
rect -1309 -617 -1297 -583
rect -1389 -623 -1297 -617
rect -1231 -583 -1139 -577
rect -1231 -617 -1219 -583
rect -1151 -617 -1139 -583
rect -1231 -623 -1139 -617
rect -1073 -583 -981 -577
rect -1073 -617 -1061 -583
rect -993 -617 -981 -583
rect -1073 -623 -981 -617
rect -915 -583 -823 -577
rect -915 -617 -903 -583
rect -835 -617 -823 -583
rect -915 -623 -823 -617
rect -757 -583 -665 -577
rect -757 -617 -745 -583
rect -677 -617 -665 -583
rect -757 -623 -665 -617
rect -599 -583 -507 -577
rect -599 -617 -587 -583
rect -519 -617 -507 -583
rect -599 -623 -507 -617
rect -441 -583 -349 -577
rect -441 -617 -429 -583
rect -361 -617 -349 -583
rect -441 -623 -349 -617
rect -283 -583 -191 -577
rect -283 -617 -271 -583
rect -203 -617 -191 -583
rect -283 -623 -191 -617
rect -125 -583 -33 -577
rect -125 -617 -113 -583
rect -45 -617 -33 -583
rect -125 -623 -33 -617
rect 33 -583 125 -577
rect 33 -617 45 -583
rect 113 -617 125 -583
rect 33 -623 125 -617
rect 191 -583 283 -577
rect 191 -617 203 -583
rect 271 -617 283 -583
rect 191 -623 283 -617
rect 349 -583 441 -577
rect 349 -617 361 -583
rect 429 -617 441 -583
rect 349 -623 441 -617
rect 507 -583 599 -577
rect 507 -617 519 -583
rect 587 -617 599 -583
rect 507 -623 599 -617
rect 665 -583 757 -577
rect 665 -617 677 -583
rect 745 -617 757 -583
rect 665 -623 757 -617
rect 823 -583 915 -577
rect 823 -617 835 -583
rect 903 -617 915 -583
rect 823 -623 915 -617
rect 981 -583 1073 -577
rect 981 -617 993 -583
rect 1061 -617 1073 -583
rect 981 -623 1073 -617
rect 1139 -583 1231 -577
rect 1139 -617 1151 -583
rect 1219 -617 1231 -583
rect 1139 -623 1231 -617
rect 1297 -583 1389 -577
rect 1297 -617 1309 -583
rect 1377 -617 1389 -583
rect 1297 -623 1389 -617
rect 1455 -583 1547 -577
rect 1455 -617 1467 -583
rect 1535 -617 1547 -583
rect 1455 -623 1547 -617
rect 1613 -583 1705 -577
rect 1613 -617 1625 -583
rect 1693 -617 1705 -583
rect 1613 -623 1705 -617
rect 1771 -583 1863 -577
rect 1771 -617 1783 -583
rect 1851 -617 1863 -583
rect 1771 -623 1863 -617
rect 1929 -583 2021 -577
rect 1929 -617 1941 -583
rect 2009 -617 2021 -583
rect 1929 -623 2021 -617
rect 2087 -583 2179 -577
rect 2087 -617 2099 -583
rect 2167 -617 2179 -583
rect 2087 -623 2179 -617
rect 2245 -583 2337 -577
rect 2245 -617 2257 -583
rect 2325 -617 2337 -583
rect 2245 -623 2337 -617
rect 2403 -583 2495 -577
rect 2403 -617 2415 -583
rect 2483 -617 2495 -583
rect 2403 -623 2495 -617
rect 2561 -583 2653 -577
rect 2561 -617 2573 -583
rect 2641 -617 2653 -583
rect 2561 -623 2653 -617
rect 2719 -583 2811 -577
rect 2719 -617 2731 -583
rect 2799 -617 2811 -583
rect 2719 -623 2811 -617
rect 2877 -583 2969 -577
rect 2877 -617 2889 -583
rect 2957 -617 2969 -583
rect 2877 -623 2969 -617
rect 3035 -583 3127 -577
rect 3035 -617 3047 -583
rect 3115 -617 3127 -583
rect 3035 -623 3127 -617
rect 3193 -583 3285 -577
rect 3193 -617 3205 -583
rect 3273 -617 3285 -583
rect 3193 -623 3285 -617
rect 3351 -583 3443 -577
rect 3351 -617 3363 -583
rect 3431 -617 3443 -583
rect 3351 -623 3443 -617
rect 3509 -583 3601 -577
rect 3509 -617 3521 -583
rect 3589 -617 3601 -583
rect 3509 -623 3601 -617
rect 3667 -583 3759 -577
rect 3667 -617 3679 -583
rect 3747 -617 3759 -583
rect 3667 -623 3759 -617
rect 3825 -583 3917 -577
rect 3825 -617 3837 -583
rect 3905 -617 3917 -583
rect 3825 -623 3917 -617
rect 3983 -583 4075 -577
rect 3983 -617 3995 -583
rect 4063 -617 4075 -583
rect 3983 -623 4075 -617
rect 4141 -583 4233 -577
rect 4141 -617 4153 -583
rect 4221 -617 4233 -583
rect 4141 -623 4233 -617
rect 4299 -583 4391 -577
rect 4299 -617 4311 -583
rect 4379 -617 4391 -583
rect 4299 -623 4391 -617
rect -4391 -691 -4299 -685
rect -4391 -725 -4379 -691
rect -4311 -725 -4299 -691
rect -4391 -731 -4299 -725
rect -4233 -691 -4141 -685
rect -4233 -725 -4221 -691
rect -4153 -725 -4141 -691
rect -4233 -731 -4141 -725
rect -4075 -691 -3983 -685
rect -4075 -725 -4063 -691
rect -3995 -725 -3983 -691
rect -4075 -731 -3983 -725
rect -3917 -691 -3825 -685
rect -3917 -725 -3905 -691
rect -3837 -725 -3825 -691
rect -3917 -731 -3825 -725
rect -3759 -691 -3667 -685
rect -3759 -725 -3747 -691
rect -3679 -725 -3667 -691
rect -3759 -731 -3667 -725
rect -3601 -691 -3509 -685
rect -3601 -725 -3589 -691
rect -3521 -725 -3509 -691
rect -3601 -731 -3509 -725
rect -3443 -691 -3351 -685
rect -3443 -725 -3431 -691
rect -3363 -725 -3351 -691
rect -3443 -731 -3351 -725
rect -3285 -691 -3193 -685
rect -3285 -725 -3273 -691
rect -3205 -725 -3193 -691
rect -3285 -731 -3193 -725
rect -3127 -691 -3035 -685
rect -3127 -725 -3115 -691
rect -3047 -725 -3035 -691
rect -3127 -731 -3035 -725
rect -2969 -691 -2877 -685
rect -2969 -725 -2957 -691
rect -2889 -725 -2877 -691
rect -2969 -731 -2877 -725
rect -2811 -691 -2719 -685
rect -2811 -725 -2799 -691
rect -2731 -725 -2719 -691
rect -2811 -731 -2719 -725
rect -2653 -691 -2561 -685
rect -2653 -725 -2641 -691
rect -2573 -725 -2561 -691
rect -2653 -731 -2561 -725
rect -2495 -691 -2403 -685
rect -2495 -725 -2483 -691
rect -2415 -725 -2403 -691
rect -2495 -731 -2403 -725
rect -2337 -691 -2245 -685
rect -2337 -725 -2325 -691
rect -2257 -725 -2245 -691
rect -2337 -731 -2245 -725
rect -2179 -691 -2087 -685
rect -2179 -725 -2167 -691
rect -2099 -725 -2087 -691
rect -2179 -731 -2087 -725
rect -2021 -691 -1929 -685
rect -2021 -725 -2009 -691
rect -1941 -725 -1929 -691
rect -2021 -731 -1929 -725
rect -1863 -691 -1771 -685
rect -1863 -725 -1851 -691
rect -1783 -725 -1771 -691
rect -1863 -731 -1771 -725
rect -1705 -691 -1613 -685
rect -1705 -725 -1693 -691
rect -1625 -725 -1613 -691
rect -1705 -731 -1613 -725
rect -1547 -691 -1455 -685
rect -1547 -725 -1535 -691
rect -1467 -725 -1455 -691
rect -1547 -731 -1455 -725
rect -1389 -691 -1297 -685
rect -1389 -725 -1377 -691
rect -1309 -725 -1297 -691
rect -1389 -731 -1297 -725
rect -1231 -691 -1139 -685
rect -1231 -725 -1219 -691
rect -1151 -725 -1139 -691
rect -1231 -731 -1139 -725
rect -1073 -691 -981 -685
rect -1073 -725 -1061 -691
rect -993 -725 -981 -691
rect -1073 -731 -981 -725
rect -915 -691 -823 -685
rect -915 -725 -903 -691
rect -835 -725 -823 -691
rect -915 -731 -823 -725
rect -757 -691 -665 -685
rect -757 -725 -745 -691
rect -677 -725 -665 -691
rect -757 -731 -665 -725
rect -599 -691 -507 -685
rect -599 -725 -587 -691
rect -519 -725 -507 -691
rect -599 -731 -507 -725
rect -441 -691 -349 -685
rect -441 -725 -429 -691
rect -361 -725 -349 -691
rect -441 -731 -349 -725
rect -283 -691 -191 -685
rect -283 -725 -271 -691
rect -203 -725 -191 -691
rect -283 -731 -191 -725
rect -125 -691 -33 -685
rect -125 -725 -113 -691
rect -45 -725 -33 -691
rect -125 -731 -33 -725
rect 33 -691 125 -685
rect 33 -725 45 -691
rect 113 -725 125 -691
rect 33 -731 125 -725
rect 191 -691 283 -685
rect 191 -725 203 -691
rect 271 -725 283 -691
rect 191 -731 283 -725
rect 349 -691 441 -685
rect 349 -725 361 -691
rect 429 -725 441 -691
rect 349 -731 441 -725
rect 507 -691 599 -685
rect 507 -725 519 -691
rect 587 -725 599 -691
rect 507 -731 599 -725
rect 665 -691 757 -685
rect 665 -725 677 -691
rect 745 -725 757 -691
rect 665 -731 757 -725
rect 823 -691 915 -685
rect 823 -725 835 -691
rect 903 -725 915 -691
rect 823 -731 915 -725
rect 981 -691 1073 -685
rect 981 -725 993 -691
rect 1061 -725 1073 -691
rect 981 -731 1073 -725
rect 1139 -691 1231 -685
rect 1139 -725 1151 -691
rect 1219 -725 1231 -691
rect 1139 -731 1231 -725
rect 1297 -691 1389 -685
rect 1297 -725 1309 -691
rect 1377 -725 1389 -691
rect 1297 -731 1389 -725
rect 1455 -691 1547 -685
rect 1455 -725 1467 -691
rect 1535 -725 1547 -691
rect 1455 -731 1547 -725
rect 1613 -691 1705 -685
rect 1613 -725 1625 -691
rect 1693 -725 1705 -691
rect 1613 -731 1705 -725
rect 1771 -691 1863 -685
rect 1771 -725 1783 -691
rect 1851 -725 1863 -691
rect 1771 -731 1863 -725
rect 1929 -691 2021 -685
rect 1929 -725 1941 -691
rect 2009 -725 2021 -691
rect 1929 -731 2021 -725
rect 2087 -691 2179 -685
rect 2087 -725 2099 -691
rect 2167 -725 2179 -691
rect 2087 -731 2179 -725
rect 2245 -691 2337 -685
rect 2245 -725 2257 -691
rect 2325 -725 2337 -691
rect 2245 -731 2337 -725
rect 2403 -691 2495 -685
rect 2403 -725 2415 -691
rect 2483 -725 2495 -691
rect 2403 -731 2495 -725
rect 2561 -691 2653 -685
rect 2561 -725 2573 -691
rect 2641 -725 2653 -691
rect 2561 -731 2653 -725
rect 2719 -691 2811 -685
rect 2719 -725 2731 -691
rect 2799 -725 2811 -691
rect 2719 -731 2811 -725
rect 2877 -691 2969 -685
rect 2877 -725 2889 -691
rect 2957 -725 2969 -691
rect 2877 -731 2969 -725
rect 3035 -691 3127 -685
rect 3035 -725 3047 -691
rect 3115 -725 3127 -691
rect 3035 -731 3127 -725
rect 3193 -691 3285 -685
rect 3193 -725 3205 -691
rect 3273 -725 3285 -691
rect 3193 -731 3285 -725
rect 3351 -691 3443 -685
rect 3351 -725 3363 -691
rect 3431 -725 3443 -691
rect 3351 -731 3443 -725
rect 3509 -691 3601 -685
rect 3509 -725 3521 -691
rect 3589 -725 3601 -691
rect 3509 -731 3601 -725
rect 3667 -691 3759 -685
rect 3667 -725 3679 -691
rect 3747 -725 3759 -691
rect 3667 -731 3759 -725
rect 3825 -691 3917 -685
rect 3825 -725 3837 -691
rect 3905 -725 3917 -691
rect 3825 -731 3917 -725
rect 3983 -691 4075 -685
rect 3983 -725 3995 -691
rect 4063 -725 4075 -691
rect 3983 -731 4075 -725
rect 4141 -691 4233 -685
rect 4141 -725 4153 -691
rect 4221 -725 4233 -691
rect 4141 -731 4233 -725
rect 4299 -691 4391 -685
rect 4299 -725 4311 -691
rect 4379 -725 4391 -691
rect 4299 -731 4391 -725
rect -4447 -784 -4401 -772
rect -4447 -960 -4441 -784
rect -4407 -960 -4401 -784
rect -4447 -972 -4401 -960
rect -4289 -784 -4243 -772
rect -4289 -960 -4283 -784
rect -4249 -960 -4243 -784
rect -4289 -972 -4243 -960
rect -4131 -784 -4085 -772
rect -4131 -960 -4125 -784
rect -4091 -960 -4085 -784
rect -4131 -972 -4085 -960
rect -3973 -784 -3927 -772
rect -3973 -960 -3967 -784
rect -3933 -960 -3927 -784
rect -3973 -972 -3927 -960
rect -3815 -784 -3769 -772
rect -3815 -960 -3809 -784
rect -3775 -960 -3769 -784
rect -3815 -972 -3769 -960
rect -3657 -784 -3611 -772
rect -3657 -960 -3651 -784
rect -3617 -960 -3611 -784
rect -3657 -972 -3611 -960
rect -3499 -784 -3453 -772
rect -3499 -960 -3493 -784
rect -3459 -960 -3453 -784
rect -3499 -972 -3453 -960
rect -3341 -784 -3295 -772
rect -3341 -960 -3335 -784
rect -3301 -960 -3295 -784
rect -3341 -972 -3295 -960
rect -3183 -784 -3137 -772
rect -3183 -960 -3177 -784
rect -3143 -960 -3137 -784
rect -3183 -972 -3137 -960
rect -3025 -784 -2979 -772
rect -3025 -960 -3019 -784
rect -2985 -960 -2979 -784
rect -3025 -972 -2979 -960
rect -2867 -784 -2821 -772
rect -2867 -960 -2861 -784
rect -2827 -960 -2821 -784
rect -2867 -972 -2821 -960
rect -2709 -784 -2663 -772
rect -2709 -960 -2703 -784
rect -2669 -960 -2663 -784
rect -2709 -972 -2663 -960
rect -2551 -784 -2505 -772
rect -2551 -960 -2545 -784
rect -2511 -960 -2505 -784
rect -2551 -972 -2505 -960
rect -2393 -784 -2347 -772
rect -2393 -960 -2387 -784
rect -2353 -960 -2347 -784
rect -2393 -972 -2347 -960
rect -2235 -784 -2189 -772
rect -2235 -960 -2229 -784
rect -2195 -960 -2189 -784
rect -2235 -972 -2189 -960
rect -2077 -784 -2031 -772
rect -2077 -960 -2071 -784
rect -2037 -960 -2031 -784
rect -2077 -972 -2031 -960
rect -1919 -784 -1873 -772
rect -1919 -960 -1913 -784
rect -1879 -960 -1873 -784
rect -1919 -972 -1873 -960
rect -1761 -784 -1715 -772
rect -1761 -960 -1755 -784
rect -1721 -960 -1715 -784
rect -1761 -972 -1715 -960
rect -1603 -784 -1557 -772
rect -1603 -960 -1597 -784
rect -1563 -960 -1557 -784
rect -1603 -972 -1557 -960
rect -1445 -784 -1399 -772
rect -1445 -960 -1439 -784
rect -1405 -960 -1399 -784
rect -1445 -972 -1399 -960
rect -1287 -784 -1241 -772
rect -1287 -960 -1281 -784
rect -1247 -960 -1241 -784
rect -1287 -972 -1241 -960
rect -1129 -784 -1083 -772
rect -1129 -960 -1123 -784
rect -1089 -960 -1083 -784
rect -1129 -972 -1083 -960
rect -971 -784 -925 -772
rect -971 -960 -965 -784
rect -931 -960 -925 -784
rect -971 -972 -925 -960
rect -813 -784 -767 -772
rect -813 -960 -807 -784
rect -773 -960 -767 -784
rect -813 -972 -767 -960
rect -655 -784 -609 -772
rect -655 -960 -649 -784
rect -615 -960 -609 -784
rect -655 -972 -609 -960
rect -497 -784 -451 -772
rect -497 -960 -491 -784
rect -457 -960 -451 -784
rect -497 -972 -451 -960
rect -339 -784 -293 -772
rect -339 -960 -333 -784
rect -299 -960 -293 -784
rect -339 -972 -293 -960
rect -181 -784 -135 -772
rect -181 -960 -175 -784
rect -141 -960 -135 -784
rect -181 -972 -135 -960
rect -23 -784 23 -772
rect -23 -960 -17 -784
rect 17 -960 23 -784
rect -23 -972 23 -960
rect 135 -784 181 -772
rect 135 -960 141 -784
rect 175 -960 181 -784
rect 135 -972 181 -960
rect 293 -784 339 -772
rect 293 -960 299 -784
rect 333 -960 339 -784
rect 293 -972 339 -960
rect 451 -784 497 -772
rect 451 -960 457 -784
rect 491 -960 497 -784
rect 451 -972 497 -960
rect 609 -784 655 -772
rect 609 -960 615 -784
rect 649 -960 655 -784
rect 609 -972 655 -960
rect 767 -784 813 -772
rect 767 -960 773 -784
rect 807 -960 813 -784
rect 767 -972 813 -960
rect 925 -784 971 -772
rect 925 -960 931 -784
rect 965 -960 971 -784
rect 925 -972 971 -960
rect 1083 -784 1129 -772
rect 1083 -960 1089 -784
rect 1123 -960 1129 -784
rect 1083 -972 1129 -960
rect 1241 -784 1287 -772
rect 1241 -960 1247 -784
rect 1281 -960 1287 -784
rect 1241 -972 1287 -960
rect 1399 -784 1445 -772
rect 1399 -960 1405 -784
rect 1439 -960 1445 -784
rect 1399 -972 1445 -960
rect 1557 -784 1603 -772
rect 1557 -960 1563 -784
rect 1597 -960 1603 -784
rect 1557 -972 1603 -960
rect 1715 -784 1761 -772
rect 1715 -960 1721 -784
rect 1755 -960 1761 -784
rect 1715 -972 1761 -960
rect 1873 -784 1919 -772
rect 1873 -960 1879 -784
rect 1913 -960 1919 -784
rect 1873 -972 1919 -960
rect 2031 -784 2077 -772
rect 2031 -960 2037 -784
rect 2071 -960 2077 -784
rect 2031 -972 2077 -960
rect 2189 -784 2235 -772
rect 2189 -960 2195 -784
rect 2229 -960 2235 -784
rect 2189 -972 2235 -960
rect 2347 -784 2393 -772
rect 2347 -960 2353 -784
rect 2387 -960 2393 -784
rect 2347 -972 2393 -960
rect 2505 -784 2551 -772
rect 2505 -960 2511 -784
rect 2545 -960 2551 -784
rect 2505 -972 2551 -960
rect 2663 -784 2709 -772
rect 2663 -960 2669 -784
rect 2703 -960 2709 -784
rect 2663 -972 2709 -960
rect 2821 -784 2867 -772
rect 2821 -960 2827 -784
rect 2861 -960 2867 -784
rect 2821 -972 2867 -960
rect 2979 -784 3025 -772
rect 2979 -960 2985 -784
rect 3019 -960 3025 -784
rect 2979 -972 3025 -960
rect 3137 -784 3183 -772
rect 3137 -960 3143 -784
rect 3177 -960 3183 -784
rect 3137 -972 3183 -960
rect 3295 -784 3341 -772
rect 3295 -960 3301 -784
rect 3335 -960 3341 -784
rect 3295 -972 3341 -960
rect 3453 -784 3499 -772
rect 3453 -960 3459 -784
rect 3493 -960 3499 -784
rect 3453 -972 3499 -960
rect 3611 -784 3657 -772
rect 3611 -960 3617 -784
rect 3651 -960 3657 -784
rect 3611 -972 3657 -960
rect 3769 -784 3815 -772
rect 3769 -960 3775 -784
rect 3809 -960 3815 -784
rect 3769 -972 3815 -960
rect 3927 -784 3973 -772
rect 3927 -960 3933 -784
rect 3967 -960 3973 -784
rect 3927 -972 3973 -960
rect 4085 -784 4131 -772
rect 4085 -960 4091 -784
rect 4125 -960 4131 -784
rect 4085 -972 4131 -960
rect 4243 -784 4289 -772
rect 4243 -960 4249 -784
rect 4283 -960 4289 -784
rect 4243 -972 4289 -960
rect 4401 -784 4447 -772
rect 4401 -960 4407 -784
rect 4441 -960 4447 -784
rect 4401 -972 4447 -960
rect -4391 -1019 -4299 -1013
rect -4391 -1053 -4379 -1019
rect -4311 -1053 -4299 -1019
rect -4391 -1059 -4299 -1053
rect -4233 -1019 -4141 -1013
rect -4233 -1053 -4221 -1019
rect -4153 -1053 -4141 -1019
rect -4233 -1059 -4141 -1053
rect -4075 -1019 -3983 -1013
rect -4075 -1053 -4063 -1019
rect -3995 -1053 -3983 -1019
rect -4075 -1059 -3983 -1053
rect -3917 -1019 -3825 -1013
rect -3917 -1053 -3905 -1019
rect -3837 -1053 -3825 -1019
rect -3917 -1059 -3825 -1053
rect -3759 -1019 -3667 -1013
rect -3759 -1053 -3747 -1019
rect -3679 -1053 -3667 -1019
rect -3759 -1059 -3667 -1053
rect -3601 -1019 -3509 -1013
rect -3601 -1053 -3589 -1019
rect -3521 -1053 -3509 -1019
rect -3601 -1059 -3509 -1053
rect -3443 -1019 -3351 -1013
rect -3443 -1053 -3431 -1019
rect -3363 -1053 -3351 -1019
rect -3443 -1059 -3351 -1053
rect -3285 -1019 -3193 -1013
rect -3285 -1053 -3273 -1019
rect -3205 -1053 -3193 -1019
rect -3285 -1059 -3193 -1053
rect -3127 -1019 -3035 -1013
rect -3127 -1053 -3115 -1019
rect -3047 -1053 -3035 -1019
rect -3127 -1059 -3035 -1053
rect -2969 -1019 -2877 -1013
rect -2969 -1053 -2957 -1019
rect -2889 -1053 -2877 -1019
rect -2969 -1059 -2877 -1053
rect -2811 -1019 -2719 -1013
rect -2811 -1053 -2799 -1019
rect -2731 -1053 -2719 -1019
rect -2811 -1059 -2719 -1053
rect -2653 -1019 -2561 -1013
rect -2653 -1053 -2641 -1019
rect -2573 -1053 -2561 -1019
rect -2653 -1059 -2561 -1053
rect -2495 -1019 -2403 -1013
rect -2495 -1053 -2483 -1019
rect -2415 -1053 -2403 -1019
rect -2495 -1059 -2403 -1053
rect -2337 -1019 -2245 -1013
rect -2337 -1053 -2325 -1019
rect -2257 -1053 -2245 -1019
rect -2337 -1059 -2245 -1053
rect -2179 -1019 -2087 -1013
rect -2179 -1053 -2167 -1019
rect -2099 -1053 -2087 -1019
rect -2179 -1059 -2087 -1053
rect -2021 -1019 -1929 -1013
rect -2021 -1053 -2009 -1019
rect -1941 -1053 -1929 -1019
rect -2021 -1059 -1929 -1053
rect -1863 -1019 -1771 -1013
rect -1863 -1053 -1851 -1019
rect -1783 -1053 -1771 -1019
rect -1863 -1059 -1771 -1053
rect -1705 -1019 -1613 -1013
rect -1705 -1053 -1693 -1019
rect -1625 -1053 -1613 -1019
rect -1705 -1059 -1613 -1053
rect -1547 -1019 -1455 -1013
rect -1547 -1053 -1535 -1019
rect -1467 -1053 -1455 -1019
rect -1547 -1059 -1455 -1053
rect -1389 -1019 -1297 -1013
rect -1389 -1053 -1377 -1019
rect -1309 -1053 -1297 -1019
rect -1389 -1059 -1297 -1053
rect -1231 -1019 -1139 -1013
rect -1231 -1053 -1219 -1019
rect -1151 -1053 -1139 -1019
rect -1231 -1059 -1139 -1053
rect -1073 -1019 -981 -1013
rect -1073 -1053 -1061 -1019
rect -993 -1053 -981 -1019
rect -1073 -1059 -981 -1053
rect -915 -1019 -823 -1013
rect -915 -1053 -903 -1019
rect -835 -1053 -823 -1019
rect -915 -1059 -823 -1053
rect -757 -1019 -665 -1013
rect -757 -1053 -745 -1019
rect -677 -1053 -665 -1019
rect -757 -1059 -665 -1053
rect -599 -1019 -507 -1013
rect -599 -1053 -587 -1019
rect -519 -1053 -507 -1019
rect -599 -1059 -507 -1053
rect -441 -1019 -349 -1013
rect -441 -1053 -429 -1019
rect -361 -1053 -349 -1019
rect -441 -1059 -349 -1053
rect -283 -1019 -191 -1013
rect -283 -1053 -271 -1019
rect -203 -1053 -191 -1019
rect -283 -1059 -191 -1053
rect -125 -1019 -33 -1013
rect -125 -1053 -113 -1019
rect -45 -1053 -33 -1019
rect -125 -1059 -33 -1053
rect 33 -1019 125 -1013
rect 33 -1053 45 -1019
rect 113 -1053 125 -1019
rect 33 -1059 125 -1053
rect 191 -1019 283 -1013
rect 191 -1053 203 -1019
rect 271 -1053 283 -1019
rect 191 -1059 283 -1053
rect 349 -1019 441 -1013
rect 349 -1053 361 -1019
rect 429 -1053 441 -1019
rect 349 -1059 441 -1053
rect 507 -1019 599 -1013
rect 507 -1053 519 -1019
rect 587 -1053 599 -1019
rect 507 -1059 599 -1053
rect 665 -1019 757 -1013
rect 665 -1053 677 -1019
rect 745 -1053 757 -1019
rect 665 -1059 757 -1053
rect 823 -1019 915 -1013
rect 823 -1053 835 -1019
rect 903 -1053 915 -1019
rect 823 -1059 915 -1053
rect 981 -1019 1073 -1013
rect 981 -1053 993 -1019
rect 1061 -1053 1073 -1019
rect 981 -1059 1073 -1053
rect 1139 -1019 1231 -1013
rect 1139 -1053 1151 -1019
rect 1219 -1053 1231 -1019
rect 1139 -1059 1231 -1053
rect 1297 -1019 1389 -1013
rect 1297 -1053 1309 -1019
rect 1377 -1053 1389 -1019
rect 1297 -1059 1389 -1053
rect 1455 -1019 1547 -1013
rect 1455 -1053 1467 -1019
rect 1535 -1053 1547 -1019
rect 1455 -1059 1547 -1053
rect 1613 -1019 1705 -1013
rect 1613 -1053 1625 -1019
rect 1693 -1053 1705 -1019
rect 1613 -1059 1705 -1053
rect 1771 -1019 1863 -1013
rect 1771 -1053 1783 -1019
rect 1851 -1053 1863 -1019
rect 1771 -1059 1863 -1053
rect 1929 -1019 2021 -1013
rect 1929 -1053 1941 -1019
rect 2009 -1053 2021 -1019
rect 1929 -1059 2021 -1053
rect 2087 -1019 2179 -1013
rect 2087 -1053 2099 -1019
rect 2167 -1053 2179 -1019
rect 2087 -1059 2179 -1053
rect 2245 -1019 2337 -1013
rect 2245 -1053 2257 -1019
rect 2325 -1053 2337 -1019
rect 2245 -1059 2337 -1053
rect 2403 -1019 2495 -1013
rect 2403 -1053 2415 -1019
rect 2483 -1053 2495 -1019
rect 2403 -1059 2495 -1053
rect 2561 -1019 2653 -1013
rect 2561 -1053 2573 -1019
rect 2641 -1053 2653 -1019
rect 2561 -1059 2653 -1053
rect 2719 -1019 2811 -1013
rect 2719 -1053 2731 -1019
rect 2799 -1053 2811 -1019
rect 2719 -1059 2811 -1053
rect 2877 -1019 2969 -1013
rect 2877 -1053 2889 -1019
rect 2957 -1053 2969 -1019
rect 2877 -1059 2969 -1053
rect 3035 -1019 3127 -1013
rect 3035 -1053 3047 -1019
rect 3115 -1053 3127 -1019
rect 3035 -1059 3127 -1053
rect 3193 -1019 3285 -1013
rect 3193 -1053 3205 -1019
rect 3273 -1053 3285 -1019
rect 3193 -1059 3285 -1053
rect 3351 -1019 3443 -1013
rect 3351 -1053 3363 -1019
rect 3431 -1053 3443 -1019
rect 3351 -1059 3443 -1053
rect 3509 -1019 3601 -1013
rect 3509 -1053 3521 -1019
rect 3589 -1053 3601 -1019
rect 3509 -1059 3601 -1053
rect 3667 -1019 3759 -1013
rect 3667 -1053 3679 -1019
rect 3747 -1053 3759 -1019
rect 3667 -1059 3759 -1053
rect 3825 -1019 3917 -1013
rect 3825 -1053 3837 -1019
rect 3905 -1053 3917 -1019
rect 3825 -1059 3917 -1053
rect 3983 -1019 4075 -1013
rect 3983 -1053 3995 -1019
rect 4063 -1053 4075 -1019
rect 3983 -1059 4075 -1053
rect 4141 -1019 4233 -1013
rect 4141 -1053 4153 -1019
rect 4221 -1053 4233 -1019
rect 4141 -1059 4233 -1053
rect 4299 -1019 4391 -1013
rect 4299 -1053 4311 -1019
rect 4379 -1053 4391 -1019
rect 4299 -1059 4391 -1053
<< properties >>
string FIXED_BBOX -4558 -1174 4558 1174
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 5 nf 56 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
