magic
tech sky130A
magscale 1 2
timestamp 1651947127
<< error_p >>
rect -3514 6331 -3454 6450
rect -3434 6331 -3374 6450
rect -3638 5369 -3374 6331
rect -3514 5250 -3454 5369
rect -3434 5250 -3374 5369
rect -3318 5366 -3112 6334
rect -1792 6331 -1732 6450
rect -1712 6331 -1652 6450
rect -1916 5369 -1652 6331
rect -1792 5250 -1732 5369
rect -1712 5250 -1652 5369
rect -1596 5366 -1390 6334
rect -70 6331 -10 6450
rect 10 6331 70 6450
rect -194 5369 70 6331
rect -70 5250 -10 5369
rect 10 5250 70 5369
rect 126 5366 332 6334
rect 1652 6331 1712 6450
rect 1732 6331 1792 6450
rect 1528 5369 1792 6331
rect 1652 5250 1712 5369
rect 1732 5250 1792 5369
rect 1848 5366 2054 6334
rect 3374 6331 3434 6450
rect 3454 6331 3514 6450
rect 3250 5369 3514 6331
rect 3374 5250 3434 5369
rect 3454 5250 3514 5369
rect 3570 5366 3776 6334
rect -3514 5031 -3454 5150
rect -3434 5031 -3374 5150
rect -3638 4069 -3374 5031
rect -3514 3950 -3454 4069
rect -3434 3950 -3374 4069
rect -3318 4066 -3112 5034
rect -1792 5031 -1732 5150
rect -1712 5031 -1652 5150
rect -1916 4069 -1652 5031
rect -1792 3950 -1732 4069
rect -1712 3950 -1652 4069
rect -1596 4066 -1390 5034
rect -70 5031 -10 5150
rect 10 5031 70 5150
rect -194 4069 70 5031
rect -70 3950 -10 4069
rect 10 3950 70 4069
rect 126 4066 332 5034
rect 1652 5031 1712 5150
rect 1732 5031 1792 5150
rect 1528 4069 1792 5031
rect 1652 3950 1712 4069
rect 1732 3950 1792 4069
rect 1848 4066 2054 5034
rect 3374 5031 3434 5150
rect 3454 5031 3514 5150
rect 3250 4069 3514 5031
rect 3374 3950 3434 4069
rect 3454 3950 3514 4069
rect 3570 4066 3776 5034
rect -3514 3731 -3454 3850
rect -3434 3731 -3374 3850
rect -3638 2769 -3374 3731
rect -3514 2650 -3454 2769
rect -3434 2650 -3374 2769
rect -3318 2766 -3112 3734
rect -1792 3731 -1732 3850
rect -1712 3731 -1652 3850
rect -1916 2769 -1652 3731
rect -1792 2650 -1732 2769
rect -1712 2650 -1652 2769
rect -1596 2766 -1390 3734
rect -70 3731 -10 3850
rect 10 3731 70 3850
rect -194 2769 70 3731
rect -70 2650 -10 2769
rect 10 2650 70 2769
rect 126 2766 332 3734
rect 1652 3731 1712 3850
rect 1732 3731 1792 3850
rect 1528 2769 1792 3731
rect 1652 2650 1712 2769
rect 1732 2650 1792 2769
rect 1848 2766 2054 3734
rect 3374 3731 3434 3850
rect 3454 3731 3514 3850
rect 3250 2769 3514 3731
rect 3374 2650 3434 2769
rect 3454 2650 3514 2769
rect 3570 2766 3776 3734
rect -3514 2431 -3454 2550
rect -3434 2431 -3374 2550
rect -3638 1469 -3374 2431
rect -3514 1350 -3454 1469
rect -3434 1350 -3374 1469
rect -3318 1466 -3112 2434
rect -1792 2431 -1732 2550
rect -1712 2431 -1652 2550
rect -1916 1469 -1652 2431
rect -1792 1350 -1732 1469
rect -1712 1350 -1652 1469
rect -1596 1466 -1390 2434
rect -70 2431 -10 2550
rect 10 2431 70 2550
rect -194 1469 70 2431
rect -70 1350 -10 1469
rect 10 1350 70 1469
rect 126 1466 332 2434
rect 1652 2431 1712 2550
rect 1732 2431 1792 2550
rect 1528 1469 1792 2431
rect 1652 1350 1712 1469
rect 1732 1350 1792 1469
rect 1848 1466 2054 2434
rect 3374 2431 3434 2550
rect 3454 2431 3514 2550
rect 3250 1469 3514 2431
rect 3374 1350 3434 1469
rect 3454 1350 3514 1469
rect 3570 1466 3776 2434
rect -3514 1131 -3454 1250
rect -3434 1131 -3374 1250
rect -3638 169 -3374 1131
rect -3514 50 -3454 169
rect -3434 50 -3374 169
rect -3318 166 -3112 1134
rect -1792 1131 -1732 1250
rect -1712 1131 -1652 1250
rect -1916 169 -1652 1131
rect -1792 50 -1732 169
rect -1712 50 -1652 169
rect -1596 166 -1390 1134
rect -70 1131 -10 1250
rect 10 1131 70 1250
rect -194 169 70 1131
rect -70 50 -10 169
rect 10 50 70 169
rect 126 166 332 1134
rect 1652 1131 1712 1250
rect 1732 1131 1792 1250
rect 1528 169 1792 1131
rect 1652 50 1712 169
rect 1732 50 1792 169
rect 1848 166 2054 1134
rect 3374 1131 3434 1250
rect 3454 1131 3514 1250
rect 3250 169 3514 1131
rect 3374 50 3434 169
rect 3454 50 3514 169
rect 3570 166 3776 1134
rect -3514 -169 -3454 -50
rect -3434 -169 -3374 -50
rect -3638 -1131 -3374 -169
rect -3514 -1250 -3454 -1131
rect -3434 -1250 -3374 -1131
rect -3318 -1134 -3112 -166
rect -1792 -169 -1732 -50
rect -1712 -169 -1652 -50
rect -1916 -1131 -1652 -169
rect -1792 -1250 -1732 -1131
rect -1712 -1250 -1652 -1131
rect -1596 -1134 -1390 -166
rect -70 -169 -10 -50
rect 10 -169 70 -50
rect -194 -1131 70 -169
rect -70 -1250 -10 -1131
rect 10 -1250 70 -1131
rect 126 -1134 332 -166
rect 1652 -169 1712 -50
rect 1732 -169 1792 -50
rect 1528 -1131 1792 -169
rect 1652 -1250 1712 -1131
rect 1732 -1250 1792 -1131
rect 1848 -1134 2054 -166
rect 3374 -169 3434 -50
rect 3454 -169 3514 -50
rect 3250 -1131 3514 -169
rect 3374 -1250 3434 -1131
rect 3454 -1250 3514 -1131
rect 3570 -1134 3776 -166
rect -3514 -1469 -3454 -1350
rect -3434 -1469 -3374 -1350
rect -3638 -2431 -3374 -1469
rect -3514 -2550 -3454 -2431
rect -3434 -2550 -3374 -2431
rect -3318 -2434 -3112 -1466
rect -1792 -1469 -1732 -1350
rect -1712 -1469 -1652 -1350
rect -1916 -2431 -1652 -1469
rect -1792 -2550 -1732 -2431
rect -1712 -2550 -1652 -2431
rect -1596 -2434 -1390 -1466
rect -70 -1469 -10 -1350
rect 10 -1469 70 -1350
rect -194 -2431 70 -1469
rect -70 -2550 -10 -2431
rect 10 -2550 70 -2431
rect 126 -2434 332 -1466
rect 1652 -1469 1712 -1350
rect 1732 -1469 1792 -1350
rect 1528 -2431 1792 -1469
rect 1652 -2550 1712 -2431
rect 1732 -2550 1792 -2431
rect 1848 -2434 2054 -1466
rect 3374 -1469 3434 -1350
rect 3454 -1469 3514 -1350
rect 3250 -2431 3514 -1469
rect 3374 -2550 3434 -2431
rect 3454 -2550 3514 -2431
rect 3570 -2434 3776 -1466
rect -3514 -2769 -3454 -2650
rect -3434 -2769 -3374 -2650
rect -3638 -3731 -3374 -2769
rect -3514 -3850 -3454 -3731
rect -3434 -3850 -3374 -3731
rect -3318 -3734 -3112 -2766
rect -1792 -2769 -1732 -2650
rect -1712 -2769 -1652 -2650
rect -1916 -3731 -1652 -2769
rect -1792 -3850 -1732 -3731
rect -1712 -3850 -1652 -3731
rect -1596 -3734 -1390 -2766
rect -70 -2769 -10 -2650
rect 10 -2769 70 -2650
rect -194 -3731 70 -2769
rect -70 -3850 -10 -3731
rect 10 -3850 70 -3731
rect 126 -3734 332 -2766
rect 1652 -2769 1712 -2650
rect 1732 -2769 1792 -2650
rect 1528 -3731 1792 -2769
rect 1652 -3850 1712 -3731
rect 1732 -3850 1792 -3731
rect 1848 -3734 2054 -2766
rect 3374 -2769 3434 -2650
rect 3454 -2769 3514 -2650
rect 3250 -3731 3514 -2769
rect 3374 -3850 3434 -3731
rect 3454 -3850 3514 -3731
rect 3570 -3734 3776 -2766
rect -3514 -4069 -3454 -3950
rect -3434 -4069 -3374 -3950
rect -3638 -5031 -3374 -4069
rect -3514 -5150 -3454 -5031
rect -3434 -5150 -3374 -5031
rect -3318 -5034 -3112 -4066
rect -1792 -4069 -1732 -3950
rect -1712 -4069 -1652 -3950
rect -1916 -5031 -1652 -4069
rect -1792 -5150 -1732 -5031
rect -1712 -5150 -1652 -5031
rect -1596 -5034 -1390 -4066
rect -70 -4069 -10 -3950
rect 10 -4069 70 -3950
rect -194 -5031 70 -4069
rect -70 -5150 -10 -5031
rect 10 -5150 70 -5031
rect 126 -5034 332 -4066
rect 1652 -4069 1712 -3950
rect 1732 -4069 1792 -3950
rect 1528 -5031 1792 -4069
rect 1652 -5150 1712 -5031
rect 1732 -5150 1792 -5031
rect 1848 -5034 2054 -4066
rect 3374 -4069 3434 -3950
rect 3454 -4069 3514 -3950
rect 3250 -5031 3514 -4069
rect 3374 -5150 3434 -5031
rect 3454 -5150 3514 -5031
rect 3570 -5034 3776 -4066
rect -3514 -5369 -3454 -5250
rect -3434 -5369 -3374 -5250
rect -3638 -6331 -3374 -5369
rect -3514 -6450 -3454 -6331
rect -3434 -6450 -3374 -6331
rect -3318 -6334 -3112 -5366
rect -1792 -5369 -1732 -5250
rect -1712 -5369 -1652 -5250
rect -1916 -6331 -1652 -5369
rect -1792 -6450 -1732 -6331
rect -1712 -6450 -1652 -6331
rect -1596 -6334 -1390 -5366
rect -70 -5369 -10 -5250
rect 10 -5369 70 -5250
rect -194 -6331 70 -5369
rect -70 -6450 -10 -6331
rect 10 -6450 70 -6331
rect 126 -6334 332 -5366
rect 1652 -5369 1712 -5250
rect 1732 -5369 1792 -5250
rect 1528 -6331 1792 -5369
rect 1652 -6450 1712 -6331
rect 1732 -6450 1792 -6331
rect 1848 -6334 2054 -5366
rect 3374 -5369 3434 -5250
rect 3454 -5369 3514 -5250
rect 3250 -6331 3514 -5369
rect 3374 -6450 3434 -6331
rect 3454 -6450 3514 -6331
rect 3570 -6334 3776 -5366
<< metal4 >>
rect -5156 6289 -3454 6450
rect -5156 5411 -3710 6289
rect -3474 5411 -3454 6289
rect -5156 5250 -3454 5411
rect -3434 6289 -1732 6450
rect -3434 5411 -1988 6289
rect -1752 5411 -1732 6289
rect -3434 5250 -1732 5411
rect -1712 6289 -10 6450
rect -1712 5411 -266 6289
rect -30 5411 -10 6289
rect -1712 5250 -10 5411
rect 10 6289 1712 6450
rect 10 5411 1456 6289
rect 1692 5411 1712 6289
rect 10 5250 1712 5411
rect 1732 6289 3434 6450
rect 1732 5411 3178 6289
rect 3414 5411 3434 6289
rect 1732 5250 3434 5411
rect 3454 6289 5156 6450
rect 3454 5411 4900 6289
rect 5136 5411 5156 6289
rect 3454 5250 5156 5411
rect -5156 4989 -3454 5150
rect -5156 4111 -3710 4989
rect -3474 4111 -3454 4989
rect -5156 3950 -3454 4111
rect -3434 4989 -1732 5150
rect -3434 4111 -1988 4989
rect -1752 4111 -1732 4989
rect -3434 3950 -1732 4111
rect -1712 4989 -10 5150
rect -1712 4111 -266 4989
rect -30 4111 -10 4989
rect -1712 3950 -10 4111
rect 10 4989 1712 5150
rect 10 4111 1456 4989
rect 1692 4111 1712 4989
rect 10 3950 1712 4111
rect 1732 4989 3434 5150
rect 1732 4111 3178 4989
rect 3414 4111 3434 4989
rect 1732 3950 3434 4111
rect 3454 4989 5156 5150
rect 3454 4111 4900 4989
rect 5136 4111 5156 4989
rect 3454 3950 5156 4111
rect -5156 3689 -3454 3850
rect -5156 2811 -3710 3689
rect -3474 2811 -3454 3689
rect -5156 2650 -3454 2811
rect -3434 3689 -1732 3850
rect -3434 2811 -1988 3689
rect -1752 2811 -1732 3689
rect -3434 2650 -1732 2811
rect -1712 3689 -10 3850
rect -1712 2811 -266 3689
rect -30 2811 -10 3689
rect -1712 2650 -10 2811
rect 10 3689 1712 3850
rect 10 2811 1456 3689
rect 1692 2811 1712 3689
rect 10 2650 1712 2811
rect 1732 3689 3434 3850
rect 1732 2811 3178 3689
rect 3414 2811 3434 3689
rect 1732 2650 3434 2811
rect 3454 3689 5156 3850
rect 3454 2811 4900 3689
rect 5136 2811 5156 3689
rect 3454 2650 5156 2811
rect -5156 2389 -3454 2550
rect -5156 1511 -3710 2389
rect -3474 1511 -3454 2389
rect -5156 1350 -3454 1511
rect -3434 2389 -1732 2550
rect -3434 1511 -1988 2389
rect -1752 1511 -1732 2389
rect -3434 1350 -1732 1511
rect -1712 2389 -10 2550
rect -1712 1511 -266 2389
rect -30 1511 -10 2389
rect -1712 1350 -10 1511
rect 10 2389 1712 2550
rect 10 1511 1456 2389
rect 1692 1511 1712 2389
rect 10 1350 1712 1511
rect 1732 2389 3434 2550
rect 1732 1511 3178 2389
rect 3414 1511 3434 2389
rect 1732 1350 3434 1511
rect 3454 2389 5156 2550
rect 3454 1511 4900 2389
rect 5136 1511 5156 2389
rect 3454 1350 5156 1511
rect -5156 1089 -3454 1250
rect -5156 211 -3710 1089
rect -3474 211 -3454 1089
rect -5156 50 -3454 211
rect -3434 1089 -1732 1250
rect -3434 211 -1988 1089
rect -1752 211 -1732 1089
rect -3434 50 -1732 211
rect -1712 1089 -10 1250
rect -1712 211 -266 1089
rect -30 211 -10 1089
rect -1712 50 -10 211
rect 10 1089 1712 1250
rect 10 211 1456 1089
rect 1692 211 1712 1089
rect 10 50 1712 211
rect 1732 1089 3434 1250
rect 1732 211 3178 1089
rect 3414 211 3434 1089
rect 1732 50 3434 211
rect 3454 1089 5156 1250
rect 3454 211 4900 1089
rect 5136 211 5156 1089
rect 3454 50 5156 211
rect -5156 -211 -3454 -50
rect -5156 -1089 -3710 -211
rect -3474 -1089 -3454 -211
rect -5156 -1250 -3454 -1089
rect -3434 -211 -1732 -50
rect -3434 -1089 -1988 -211
rect -1752 -1089 -1732 -211
rect -3434 -1250 -1732 -1089
rect -1712 -211 -10 -50
rect -1712 -1089 -266 -211
rect -30 -1089 -10 -211
rect -1712 -1250 -10 -1089
rect 10 -211 1712 -50
rect 10 -1089 1456 -211
rect 1692 -1089 1712 -211
rect 10 -1250 1712 -1089
rect 1732 -211 3434 -50
rect 1732 -1089 3178 -211
rect 3414 -1089 3434 -211
rect 1732 -1250 3434 -1089
rect 3454 -211 5156 -50
rect 3454 -1089 4900 -211
rect 5136 -1089 5156 -211
rect 3454 -1250 5156 -1089
rect -5156 -1511 -3454 -1350
rect -5156 -2389 -3710 -1511
rect -3474 -2389 -3454 -1511
rect -5156 -2550 -3454 -2389
rect -3434 -1511 -1732 -1350
rect -3434 -2389 -1988 -1511
rect -1752 -2389 -1732 -1511
rect -3434 -2550 -1732 -2389
rect -1712 -1511 -10 -1350
rect -1712 -2389 -266 -1511
rect -30 -2389 -10 -1511
rect -1712 -2550 -10 -2389
rect 10 -1511 1712 -1350
rect 10 -2389 1456 -1511
rect 1692 -2389 1712 -1511
rect 10 -2550 1712 -2389
rect 1732 -1511 3434 -1350
rect 1732 -2389 3178 -1511
rect 3414 -2389 3434 -1511
rect 1732 -2550 3434 -2389
rect 3454 -1511 5156 -1350
rect 3454 -2389 4900 -1511
rect 5136 -2389 5156 -1511
rect 3454 -2550 5156 -2389
rect -5156 -2811 -3454 -2650
rect -5156 -3689 -3710 -2811
rect -3474 -3689 -3454 -2811
rect -5156 -3850 -3454 -3689
rect -3434 -2811 -1732 -2650
rect -3434 -3689 -1988 -2811
rect -1752 -3689 -1732 -2811
rect -3434 -3850 -1732 -3689
rect -1712 -2811 -10 -2650
rect -1712 -3689 -266 -2811
rect -30 -3689 -10 -2811
rect -1712 -3850 -10 -3689
rect 10 -2811 1712 -2650
rect 10 -3689 1456 -2811
rect 1692 -3689 1712 -2811
rect 10 -3850 1712 -3689
rect 1732 -2811 3434 -2650
rect 1732 -3689 3178 -2811
rect 3414 -3689 3434 -2811
rect 1732 -3850 3434 -3689
rect 3454 -2811 5156 -2650
rect 3454 -3689 4900 -2811
rect 5136 -3689 5156 -2811
rect 3454 -3850 5156 -3689
rect -5156 -4111 -3454 -3950
rect -5156 -4989 -3710 -4111
rect -3474 -4989 -3454 -4111
rect -5156 -5150 -3454 -4989
rect -3434 -4111 -1732 -3950
rect -3434 -4989 -1988 -4111
rect -1752 -4989 -1732 -4111
rect -3434 -5150 -1732 -4989
rect -1712 -4111 -10 -3950
rect -1712 -4989 -266 -4111
rect -30 -4989 -10 -4111
rect -1712 -5150 -10 -4989
rect 10 -4111 1712 -3950
rect 10 -4989 1456 -4111
rect 1692 -4989 1712 -4111
rect 10 -5150 1712 -4989
rect 1732 -4111 3434 -3950
rect 1732 -4989 3178 -4111
rect 3414 -4989 3434 -4111
rect 1732 -5150 3434 -4989
rect 3454 -4111 5156 -3950
rect 3454 -4989 4900 -4111
rect 5136 -4989 5156 -4111
rect 3454 -5150 5156 -4989
rect -5156 -5411 -3454 -5250
rect -5156 -6289 -3710 -5411
rect -3474 -6289 -3454 -5411
rect -5156 -6450 -3454 -6289
rect -3434 -5411 -1732 -5250
rect -3434 -6289 -1988 -5411
rect -1752 -6289 -1732 -5411
rect -3434 -6450 -1732 -6289
rect -1712 -5411 -10 -5250
rect -1712 -6289 -266 -5411
rect -30 -6289 -10 -5411
rect -1712 -6450 -10 -6289
rect 10 -5411 1712 -5250
rect 10 -6289 1456 -5411
rect 1692 -6289 1712 -5411
rect 10 -6450 1712 -6289
rect 1732 -5411 3434 -5250
rect 1732 -6289 3178 -5411
rect 3414 -6289 3434 -5411
rect 1732 -6450 3434 -6289
rect 3454 -5411 5156 -5250
rect 3454 -6289 4900 -5411
rect 5136 -6289 5156 -5411
rect 3454 -6450 5156 -6289
<< via4 >>
rect -3710 5411 -3474 6289
rect -1988 5411 -1752 6289
rect -266 5411 -30 6289
rect 1456 5411 1692 6289
rect 3178 5411 3414 6289
rect 4900 5411 5136 6289
rect -3710 4111 -3474 4989
rect -1988 4111 -1752 4989
rect -266 4111 -30 4989
rect 1456 4111 1692 4989
rect 3178 4111 3414 4989
rect 4900 4111 5136 4989
rect -3710 2811 -3474 3689
rect -1988 2811 -1752 3689
rect -266 2811 -30 3689
rect 1456 2811 1692 3689
rect 3178 2811 3414 3689
rect 4900 2811 5136 3689
rect -3710 1511 -3474 2389
rect -1988 1511 -1752 2389
rect -266 1511 -30 2389
rect 1456 1511 1692 2389
rect 3178 1511 3414 2389
rect 4900 1511 5136 2389
rect -3710 211 -3474 1089
rect -1988 211 -1752 1089
rect -266 211 -30 1089
rect 1456 211 1692 1089
rect 3178 211 3414 1089
rect 4900 211 5136 1089
rect -3710 -1089 -3474 -211
rect -1988 -1089 -1752 -211
rect -266 -1089 -30 -211
rect 1456 -1089 1692 -211
rect 3178 -1089 3414 -211
rect 4900 -1089 5136 -211
rect -3710 -2389 -3474 -1511
rect -1988 -2389 -1752 -1511
rect -266 -2389 -30 -1511
rect 1456 -2389 1692 -1511
rect 3178 -2389 3414 -1511
rect 4900 -2389 5136 -1511
rect -3710 -3689 -3474 -2811
rect -1988 -3689 -1752 -2811
rect -266 -3689 -30 -2811
rect 1456 -3689 1692 -2811
rect 3178 -3689 3414 -2811
rect 4900 -3689 5136 -2811
rect -3710 -4989 -3474 -4111
rect -1988 -4989 -1752 -4111
rect -266 -4989 -30 -4111
rect 1456 -4989 1692 -4111
rect 3178 -4989 3414 -4111
rect 4900 -4989 5136 -4111
rect -3710 -6289 -3474 -5411
rect -1988 -6289 -1752 -5411
rect -266 -6289 -30 -5411
rect 1456 -6289 1692 -5411
rect 3178 -6289 3414 -5411
rect 4900 -6289 5136 -5411
<< mimcap2 >>
rect -5056 6310 -4056 6350
rect -5056 5390 -5016 6310
rect -4096 5390 -4056 6310
rect -5056 5350 -4056 5390
rect -3334 6310 -2334 6350
rect -3334 5390 -3294 6310
rect -2374 5390 -2334 6310
rect -3334 5350 -2334 5390
rect -1612 6310 -612 6350
rect -1612 5390 -1572 6310
rect -652 5390 -612 6310
rect -1612 5350 -612 5390
rect 110 6310 1110 6350
rect 110 5390 150 6310
rect 1070 5390 1110 6310
rect 110 5350 1110 5390
rect 1832 6310 2832 6350
rect 1832 5390 1872 6310
rect 2792 5390 2832 6310
rect 1832 5350 2832 5390
rect 3554 6310 4554 6350
rect 3554 5390 3594 6310
rect 4514 5390 4554 6310
rect 3554 5350 4554 5390
rect -5056 5010 -4056 5050
rect -5056 4090 -5016 5010
rect -4096 4090 -4056 5010
rect -5056 4050 -4056 4090
rect -3334 5010 -2334 5050
rect -3334 4090 -3294 5010
rect -2374 4090 -2334 5010
rect -3334 4050 -2334 4090
rect -1612 5010 -612 5050
rect -1612 4090 -1572 5010
rect -652 4090 -612 5010
rect -1612 4050 -612 4090
rect 110 5010 1110 5050
rect 110 4090 150 5010
rect 1070 4090 1110 5010
rect 110 4050 1110 4090
rect 1832 5010 2832 5050
rect 1832 4090 1872 5010
rect 2792 4090 2832 5010
rect 1832 4050 2832 4090
rect 3554 5010 4554 5050
rect 3554 4090 3594 5010
rect 4514 4090 4554 5010
rect 3554 4050 4554 4090
rect -5056 3710 -4056 3750
rect -5056 2790 -5016 3710
rect -4096 2790 -4056 3710
rect -5056 2750 -4056 2790
rect -3334 3710 -2334 3750
rect -3334 2790 -3294 3710
rect -2374 2790 -2334 3710
rect -3334 2750 -2334 2790
rect -1612 3710 -612 3750
rect -1612 2790 -1572 3710
rect -652 2790 -612 3710
rect -1612 2750 -612 2790
rect 110 3710 1110 3750
rect 110 2790 150 3710
rect 1070 2790 1110 3710
rect 110 2750 1110 2790
rect 1832 3710 2832 3750
rect 1832 2790 1872 3710
rect 2792 2790 2832 3710
rect 1832 2750 2832 2790
rect 3554 3710 4554 3750
rect 3554 2790 3594 3710
rect 4514 2790 4554 3710
rect 3554 2750 4554 2790
rect -5056 2410 -4056 2450
rect -5056 1490 -5016 2410
rect -4096 1490 -4056 2410
rect -5056 1450 -4056 1490
rect -3334 2410 -2334 2450
rect -3334 1490 -3294 2410
rect -2374 1490 -2334 2410
rect -3334 1450 -2334 1490
rect -1612 2410 -612 2450
rect -1612 1490 -1572 2410
rect -652 1490 -612 2410
rect -1612 1450 -612 1490
rect 110 2410 1110 2450
rect 110 1490 150 2410
rect 1070 1490 1110 2410
rect 110 1450 1110 1490
rect 1832 2410 2832 2450
rect 1832 1490 1872 2410
rect 2792 1490 2832 2410
rect 1832 1450 2832 1490
rect 3554 2410 4554 2450
rect 3554 1490 3594 2410
rect 4514 1490 4554 2410
rect 3554 1450 4554 1490
rect -5056 1110 -4056 1150
rect -5056 190 -5016 1110
rect -4096 190 -4056 1110
rect -5056 150 -4056 190
rect -3334 1110 -2334 1150
rect -3334 190 -3294 1110
rect -2374 190 -2334 1110
rect -3334 150 -2334 190
rect -1612 1110 -612 1150
rect -1612 190 -1572 1110
rect -652 190 -612 1110
rect -1612 150 -612 190
rect 110 1110 1110 1150
rect 110 190 150 1110
rect 1070 190 1110 1110
rect 110 150 1110 190
rect 1832 1110 2832 1150
rect 1832 190 1872 1110
rect 2792 190 2832 1110
rect 1832 150 2832 190
rect 3554 1110 4554 1150
rect 3554 190 3594 1110
rect 4514 190 4554 1110
rect 3554 150 4554 190
rect -5056 -190 -4056 -150
rect -5056 -1110 -5016 -190
rect -4096 -1110 -4056 -190
rect -5056 -1150 -4056 -1110
rect -3334 -190 -2334 -150
rect -3334 -1110 -3294 -190
rect -2374 -1110 -2334 -190
rect -3334 -1150 -2334 -1110
rect -1612 -190 -612 -150
rect -1612 -1110 -1572 -190
rect -652 -1110 -612 -190
rect -1612 -1150 -612 -1110
rect 110 -190 1110 -150
rect 110 -1110 150 -190
rect 1070 -1110 1110 -190
rect 110 -1150 1110 -1110
rect 1832 -190 2832 -150
rect 1832 -1110 1872 -190
rect 2792 -1110 2832 -190
rect 1832 -1150 2832 -1110
rect 3554 -190 4554 -150
rect 3554 -1110 3594 -190
rect 4514 -1110 4554 -190
rect 3554 -1150 4554 -1110
rect -5056 -1490 -4056 -1450
rect -5056 -2410 -5016 -1490
rect -4096 -2410 -4056 -1490
rect -5056 -2450 -4056 -2410
rect -3334 -1490 -2334 -1450
rect -3334 -2410 -3294 -1490
rect -2374 -2410 -2334 -1490
rect -3334 -2450 -2334 -2410
rect -1612 -1490 -612 -1450
rect -1612 -2410 -1572 -1490
rect -652 -2410 -612 -1490
rect -1612 -2450 -612 -2410
rect 110 -1490 1110 -1450
rect 110 -2410 150 -1490
rect 1070 -2410 1110 -1490
rect 110 -2450 1110 -2410
rect 1832 -1490 2832 -1450
rect 1832 -2410 1872 -1490
rect 2792 -2410 2832 -1490
rect 1832 -2450 2832 -2410
rect 3554 -1490 4554 -1450
rect 3554 -2410 3594 -1490
rect 4514 -2410 4554 -1490
rect 3554 -2450 4554 -2410
rect -5056 -2790 -4056 -2750
rect -5056 -3710 -5016 -2790
rect -4096 -3710 -4056 -2790
rect -5056 -3750 -4056 -3710
rect -3334 -2790 -2334 -2750
rect -3334 -3710 -3294 -2790
rect -2374 -3710 -2334 -2790
rect -3334 -3750 -2334 -3710
rect -1612 -2790 -612 -2750
rect -1612 -3710 -1572 -2790
rect -652 -3710 -612 -2790
rect -1612 -3750 -612 -3710
rect 110 -2790 1110 -2750
rect 110 -3710 150 -2790
rect 1070 -3710 1110 -2790
rect 110 -3750 1110 -3710
rect 1832 -2790 2832 -2750
rect 1832 -3710 1872 -2790
rect 2792 -3710 2832 -2790
rect 1832 -3750 2832 -3710
rect 3554 -2790 4554 -2750
rect 3554 -3710 3594 -2790
rect 4514 -3710 4554 -2790
rect 3554 -3750 4554 -3710
rect -5056 -4090 -4056 -4050
rect -5056 -5010 -5016 -4090
rect -4096 -5010 -4056 -4090
rect -5056 -5050 -4056 -5010
rect -3334 -4090 -2334 -4050
rect -3334 -5010 -3294 -4090
rect -2374 -5010 -2334 -4090
rect -3334 -5050 -2334 -5010
rect -1612 -4090 -612 -4050
rect -1612 -5010 -1572 -4090
rect -652 -5010 -612 -4090
rect -1612 -5050 -612 -5010
rect 110 -4090 1110 -4050
rect 110 -5010 150 -4090
rect 1070 -5010 1110 -4090
rect 110 -5050 1110 -5010
rect 1832 -4090 2832 -4050
rect 1832 -5010 1872 -4090
rect 2792 -5010 2832 -4090
rect 1832 -5050 2832 -5010
rect 3554 -4090 4554 -4050
rect 3554 -5010 3594 -4090
rect 4514 -5010 4554 -4090
rect 3554 -5050 4554 -5010
rect -5056 -5390 -4056 -5350
rect -5056 -6310 -5016 -5390
rect -4096 -6310 -4056 -5390
rect -5056 -6350 -4056 -6310
rect -3334 -5390 -2334 -5350
rect -3334 -6310 -3294 -5390
rect -2374 -6310 -2334 -5390
rect -3334 -6350 -2334 -6310
rect -1612 -5390 -612 -5350
rect -1612 -6310 -1572 -5390
rect -652 -6310 -612 -5390
rect -1612 -6350 -612 -6310
rect 110 -5390 1110 -5350
rect 110 -6310 150 -5390
rect 1070 -6310 1110 -5390
rect 110 -6350 1110 -6310
rect 1832 -5390 2832 -5350
rect 1832 -6310 1872 -5390
rect 2792 -6310 2832 -5390
rect 1832 -6350 2832 -6310
rect 3554 -5390 4554 -5350
rect 3554 -6310 3594 -5390
rect 4514 -6310 4554 -5390
rect 3554 -6350 4554 -6310
<< mimcap2contact >>
rect -5016 5390 -4096 6310
rect -3294 5390 -2374 6310
rect -1572 5390 -652 6310
rect 150 5390 1070 6310
rect 1872 5390 2792 6310
rect 3594 5390 4514 6310
rect -5016 4090 -4096 5010
rect -3294 4090 -2374 5010
rect -1572 4090 -652 5010
rect 150 4090 1070 5010
rect 1872 4090 2792 5010
rect 3594 4090 4514 5010
rect -5016 2790 -4096 3710
rect -3294 2790 -2374 3710
rect -1572 2790 -652 3710
rect 150 2790 1070 3710
rect 1872 2790 2792 3710
rect 3594 2790 4514 3710
rect -5016 1490 -4096 2410
rect -3294 1490 -2374 2410
rect -1572 1490 -652 2410
rect 150 1490 1070 2410
rect 1872 1490 2792 2410
rect 3594 1490 4514 2410
rect -5016 190 -4096 1110
rect -3294 190 -2374 1110
rect -1572 190 -652 1110
rect 150 190 1070 1110
rect 1872 190 2792 1110
rect 3594 190 4514 1110
rect -5016 -1110 -4096 -190
rect -3294 -1110 -2374 -190
rect -1572 -1110 -652 -190
rect 150 -1110 1070 -190
rect 1872 -1110 2792 -190
rect 3594 -1110 4514 -190
rect -5016 -2410 -4096 -1490
rect -3294 -2410 -2374 -1490
rect -1572 -2410 -652 -1490
rect 150 -2410 1070 -1490
rect 1872 -2410 2792 -1490
rect 3594 -2410 4514 -1490
rect -5016 -3710 -4096 -2790
rect -3294 -3710 -2374 -2790
rect -1572 -3710 -652 -2790
rect 150 -3710 1070 -2790
rect 1872 -3710 2792 -2790
rect 3594 -3710 4514 -2790
rect -5016 -5010 -4096 -4090
rect -3294 -5010 -2374 -4090
rect -1572 -5010 -652 -4090
rect 150 -5010 1070 -4090
rect 1872 -5010 2792 -4090
rect 3594 -5010 4514 -4090
rect -5016 -6310 -4096 -5390
rect -3294 -6310 -2374 -5390
rect -1572 -6310 -652 -5390
rect 150 -6310 1070 -5390
rect 1872 -6310 2792 -5390
rect 3594 -6310 4514 -5390
<< metal5 >>
rect -4716 6334 -4396 6500
rect -2994 6334 -2674 6500
rect -1272 6334 -952 6500
rect 450 6334 770 6500
rect 2172 6334 2492 6500
rect 3894 6334 4214 6500
rect -5040 6310 -4072 6334
rect -5040 5390 -5016 6310
rect -4096 5390 -4072 6310
rect -5040 5366 -4072 5390
rect -3752 6289 -3432 6331
rect -3752 5411 -3710 6289
rect -3474 5411 -3432 6289
rect -3752 5369 -3432 5411
rect -3318 6310 -2350 6334
rect -3318 5390 -3294 6310
rect -2374 5390 -2350 6310
rect -3318 5366 -2350 5390
rect -2030 6289 -1710 6331
rect -2030 5411 -1988 6289
rect -1752 5411 -1710 6289
rect -2030 5369 -1710 5411
rect -1596 6310 -628 6334
rect -1596 5390 -1572 6310
rect -652 5390 -628 6310
rect -1596 5366 -628 5390
rect -308 6289 12 6331
rect -308 5411 -266 6289
rect -30 5411 12 6289
rect -308 5369 12 5411
rect 126 6310 1094 6334
rect 126 5390 150 6310
rect 1070 5390 1094 6310
rect 126 5366 1094 5390
rect 1414 6289 1734 6331
rect 1414 5411 1456 6289
rect 1692 5411 1734 6289
rect 1414 5369 1734 5411
rect 1848 6310 2816 6334
rect 1848 5390 1872 6310
rect 2792 5390 2816 6310
rect 1848 5366 2816 5390
rect 3136 6289 3456 6331
rect 3136 5411 3178 6289
rect 3414 5411 3456 6289
rect 3136 5369 3456 5411
rect 3570 6310 4538 6334
rect 3570 5390 3594 6310
rect 4514 5390 4538 6310
rect 3570 5366 4538 5390
rect 4858 6289 5178 6331
rect 4858 5411 4900 6289
rect 5136 5411 5178 6289
rect 4858 5369 5178 5411
rect -4716 5034 -4396 5366
rect -2994 5034 -2674 5366
rect -1272 5034 -952 5366
rect 450 5034 770 5366
rect 2172 5034 2492 5366
rect 3894 5034 4214 5366
rect -5040 5010 -4072 5034
rect -5040 4090 -5016 5010
rect -4096 4090 -4072 5010
rect -5040 4066 -4072 4090
rect -3752 4989 -3432 5031
rect -3752 4111 -3710 4989
rect -3474 4111 -3432 4989
rect -3752 4069 -3432 4111
rect -3318 5010 -2350 5034
rect -3318 4090 -3294 5010
rect -2374 4090 -2350 5010
rect -3318 4066 -2350 4090
rect -2030 4989 -1710 5031
rect -2030 4111 -1988 4989
rect -1752 4111 -1710 4989
rect -2030 4069 -1710 4111
rect -1596 5010 -628 5034
rect -1596 4090 -1572 5010
rect -652 4090 -628 5010
rect -1596 4066 -628 4090
rect -308 4989 12 5031
rect -308 4111 -266 4989
rect -30 4111 12 4989
rect -308 4069 12 4111
rect 126 5010 1094 5034
rect 126 4090 150 5010
rect 1070 4090 1094 5010
rect 126 4066 1094 4090
rect 1414 4989 1734 5031
rect 1414 4111 1456 4989
rect 1692 4111 1734 4989
rect 1414 4069 1734 4111
rect 1848 5010 2816 5034
rect 1848 4090 1872 5010
rect 2792 4090 2816 5010
rect 1848 4066 2816 4090
rect 3136 4989 3456 5031
rect 3136 4111 3178 4989
rect 3414 4111 3456 4989
rect 3136 4069 3456 4111
rect 3570 5010 4538 5034
rect 3570 4090 3594 5010
rect 4514 4090 4538 5010
rect 3570 4066 4538 4090
rect 4858 4989 5178 5031
rect 4858 4111 4900 4989
rect 5136 4111 5178 4989
rect 4858 4069 5178 4111
rect -4716 3734 -4396 4066
rect -2994 3734 -2674 4066
rect -1272 3734 -952 4066
rect 450 3734 770 4066
rect 2172 3734 2492 4066
rect 3894 3734 4214 4066
rect -5040 3710 -4072 3734
rect -5040 2790 -5016 3710
rect -4096 2790 -4072 3710
rect -5040 2766 -4072 2790
rect -3752 3689 -3432 3731
rect -3752 2811 -3710 3689
rect -3474 2811 -3432 3689
rect -3752 2769 -3432 2811
rect -3318 3710 -2350 3734
rect -3318 2790 -3294 3710
rect -2374 2790 -2350 3710
rect -3318 2766 -2350 2790
rect -2030 3689 -1710 3731
rect -2030 2811 -1988 3689
rect -1752 2811 -1710 3689
rect -2030 2769 -1710 2811
rect -1596 3710 -628 3734
rect -1596 2790 -1572 3710
rect -652 2790 -628 3710
rect -1596 2766 -628 2790
rect -308 3689 12 3731
rect -308 2811 -266 3689
rect -30 2811 12 3689
rect -308 2769 12 2811
rect 126 3710 1094 3734
rect 126 2790 150 3710
rect 1070 2790 1094 3710
rect 126 2766 1094 2790
rect 1414 3689 1734 3731
rect 1414 2811 1456 3689
rect 1692 2811 1734 3689
rect 1414 2769 1734 2811
rect 1848 3710 2816 3734
rect 1848 2790 1872 3710
rect 2792 2790 2816 3710
rect 1848 2766 2816 2790
rect 3136 3689 3456 3731
rect 3136 2811 3178 3689
rect 3414 2811 3456 3689
rect 3136 2769 3456 2811
rect 3570 3710 4538 3734
rect 3570 2790 3594 3710
rect 4514 2790 4538 3710
rect 3570 2766 4538 2790
rect 4858 3689 5178 3731
rect 4858 2811 4900 3689
rect 5136 2811 5178 3689
rect 4858 2769 5178 2811
rect -4716 2434 -4396 2766
rect -2994 2434 -2674 2766
rect -1272 2434 -952 2766
rect 450 2434 770 2766
rect 2172 2434 2492 2766
rect 3894 2434 4214 2766
rect -5040 2410 -4072 2434
rect -5040 1490 -5016 2410
rect -4096 1490 -4072 2410
rect -5040 1466 -4072 1490
rect -3752 2389 -3432 2431
rect -3752 1511 -3710 2389
rect -3474 1511 -3432 2389
rect -3752 1469 -3432 1511
rect -3318 2410 -2350 2434
rect -3318 1490 -3294 2410
rect -2374 1490 -2350 2410
rect -3318 1466 -2350 1490
rect -2030 2389 -1710 2431
rect -2030 1511 -1988 2389
rect -1752 1511 -1710 2389
rect -2030 1469 -1710 1511
rect -1596 2410 -628 2434
rect -1596 1490 -1572 2410
rect -652 1490 -628 2410
rect -1596 1466 -628 1490
rect -308 2389 12 2431
rect -308 1511 -266 2389
rect -30 1511 12 2389
rect -308 1469 12 1511
rect 126 2410 1094 2434
rect 126 1490 150 2410
rect 1070 1490 1094 2410
rect 126 1466 1094 1490
rect 1414 2389 1734 2431
rect 1414 1511 1456 2389
rect 1692 1511 1734 2389
rect 1414 1469 1734 1511
rect 1848 2410 2816 2434
rect 1848 1490 1872 2410
rect 2792 1490 2816 2410
rect 1848 1466 2816 1490
rect 3136 2389 3456 2431
rect 3136 1511 3178 2389
rect 3414 1511 3456 2389
rect 3136 1469 3456 1511
rect 3570 2410 4538 2434
rect 3570 1490 3594 2410
rect 4514 1490 4538 2410
rect 3570 1466 4538 1490
rect 4858 2389 5178 2431
rect 4858 1511 4900 2389
rect 5136 1511 5178 2389
rect 4858 1469 5178 1511
rect -4716 1134 -4396 1466
rect -2994 1134 -2674 1466
rect -1272 1134 -952 1466
rect 450 1134 770 1466
rect 2172 1134 2492 1466
rect 3894 1134 4214 1466
rect -5040 1110 -4072 1134
rect -5040 190 -5016 1110
rect -4096 190 -4072 1110
rect -5040 166 -4072 190
rect -3752 1089 -3432 1131
rect -3752 211 -3710 1089
rect -3474 211 -3432 1089
rect -3752 169 -3432 211
rect -3318 1110 -2350 1134
rect -3318 190 -3294 1110
rect -2374 190 -2350 1110
rect -3318 166 -2350 190
rect -2030 1089 -1710 1131
rect -2030 211 -1988 1089
rect -1752 211 -1710 1089
rect -2030 169 -1710 211
rect -1596 1110 -628 1134
rect -1596 190 -1572 1110
rect -652 190 -628 1110
rect -1596 166 -628 190
rect -308 1089 12 1131
rect -308 211 -266 1089
rect -30 211 12 1089
rect -308 169 12 211
rect 126 1110 1094 1134
rect 126 190 150 1110
rect 1070 190 1094 1110
rect 126 166 1094 190
rect 1414 1089 1734 1131
rect 1414 211 1456 1089
rect 1692 211 1734 1089
rect 1414 169 1734 211
rect 1848 1110 2816 1134
rect 1848 190 1872 1110
rect 2792 190 2816 1110
rect 1848 166 2816 190
rect 3136 1089 3456 1131
rect 3136 211 3178 1089
rect 3414 211 3456 1089
rect 3136 169 3456 211
rect 3570 1110 4538 1134
rect 3570 190 3594 1110
rect 4514 190 4538 1110
rect 3570 166 4538 190
rect 4858 1089 5178 1131
rect 4858 211 4900 1089
rect 5136 211 5178 1089
rect 4858 169 5178 211
rect -4716 -166 -4396 166
rect -2994 -166 -2674 166
rect -1272 -166 -952 166
rect 450 -166 770 166
rect 2172 -166 2492 166
rect 3894 -166 4214 166
rect -5040 -190 -4072 -166
rect -5040 -1110 -5016 -190
rect -4096 -1110 -4072 -190
rect -5040 -1134 -4072 -1110
rect -3752 -211 -3432 -169
rect -3752 -1089 -3710 -211
rect -3474 -1089 -3432 -211
rect -3752 -1131 -3432 -1089
rect -3318 -190 -2350 -166
rect -3318 -1110 -3294 -190
rect -2374 -1110 -2350 -190
rect -3318 -1134 -2350 -1110
rect -2030 -211 -1710 -169
rect -2030 -1089 -1988 -211
rect -1752 -1089 -1710 -211
rect -2030 -1131 -1710 -1089
rect -1596 -190 -628 -166
rect -1596 -1110 -1572 -190
rect -652 -1110 -628 -190
rect -1596 -1134 -628 -1110
rect -308 -211 12 -169
rect -308 -1089 -266 -211
rect -30 -1089 12 -211
rect -308 -1131 12 -1089
rect 126 -190 1094 -166
rect 126 -1110 150 -190
rect 1070 -1110 1094 -190
rect 126 -1134 1094 -1110
rect 1414 -211 1734 -169
rect 1414 -1089 1456 -211
rect 1692 -1089 1734 -211
rect 1414 -1131 1734 -1089
rect 1848 -190 2816 -166
rect 1848 -1110 1872 -190
rect 2792 -1110 2816 -190
rect 1848 -1134 2816 -1110
rect 3136 -211 3456 -169
rect 3136 -1089 3178 -211
rect 3414 -1089 3456 -211
rect 3136 -1131 3456 -1089
rect 3570 -190 4538 -166
rect 3570 -1110 3594 -190
rect 4514 -1110 4538 -190
rect 3570 -1134 4538 -1110
rect 4858 -211 5178 -169
rect 4858 -1089 4900 -211
rect 5136 -1089 5178 -211
rect 4858 -1131 5178 -1089
rect -4716 -1466 -4396 -1134
rect -2994 -1466 -2674 -1134
rect -1272 -1466 -952 -1134
rect 450 -1466 770 -1134
rect 2172 -1466 2492 -1134
rect 3894 -1466 4214 -1134
rect -5040 -1490 -4072 -1466
rect -5040 -2410 -5016 -1490
rect -4096 -2410 -4072 -1490
rect -5040 -2434 -4072 -2410
rect -3752 -1511 -3432 -1469
rect -3752 -2389 -3710 -1511
rect -3474 -2389 -3432 -1511
rect -3752 -2431 -3432 -2389
rect -3318 -1490 -2350 -1466
rect -3318 -2410 -3294 -1490
rect -2374 -2410 -2350 -1490
rect -3318 -2434 -2350 -2410
rect -2030 -1511 -1710 -1469
rect -2030 -2389 -1988 -1511
rect -1752 -2389 -1710 -1511
rect -2030 -2431 -1710 -2389
rect -1596 -1490 -628 -1466
rect -1596 -2410 -1572 -1490
rect -652 -2410 -628 -1490
rect -1596 -2434 -628 -2410
rect -308 -1511 12 -1469
rect -308 -2389 -266 -1511
rect -30 -2389 12 -1511
rect -308 -2431 12 -2389
rect 126 -1490 1094 -1466
rect 126 -2410 150 -1490
rect 1070 -2410 1094 -1490
rect 126 -2434 1094 -2410
rect 1414 -1511 1734 -1469
rect 1414 -2389 1456 -1511
rect 1692 -2389 1734 -1511
rect 1414 -2431 1734 -2389
rect 1848 -1490 2816 -1466
rect 1848 -2410 1872 -1490
rect 2792 -2410 2816 -1490
rect 1848 -2434 2816 -2410
rect 3136 -1511 3456 -1469
rect 3136 -2389 3178 -1511
rect 3414 -2389 3456 -1511
rect 3136 -2431 3456 -2389
rect 3570 -1490 4538 -1466
rect 3570 -2410 3594 -1490
rect 4514 -2410 4538 -1490
rect 3570 -2434 4538 -2410
rect 4858 -1511 5178 -1469
rect 4858 -2389 4900 -1511
rect 5136 -2389 5178 -1511
rect 4858 -2431 5178 -2389
rect -4716 -2766 -4396 -2434
rect -2994 -2766 -2674 -2434
rect -1272 -2766 -952 -2434
rect 450 -2766 770 -2434
rect 2172 -2766 2492 -2434
rect 3894 -2766 4214 -2434
rect -5040 -2790 -4072 -2766
rect -5040 -3710 -5016 -2790
rect -4096 -3710 -4072 -2790
rect -5040 -3734 -4072 -3710
rect -3752 -2811 -3432 -2769
rect -3752 -3689 -3710 -2811
rect -3474 -3689 -3432 -2811
rect -3752 -3731 -3432 -3689
rect -3318 -2790 -2350 -2766
rect -3318 -3710 -3294 -2790
rect -2374 -3710 -2350 -2790
rect -3318 -3734 -2350 -3710
rect -2030 -2811 -1710 -2769
rect -2030 -3689 -1988 -2811
rect -1752 -3689 -1710 -2811
rect -2030 -3731 -1710 -3689
rect -1596 -2790 -628 -2766
rect -1596 -3710 -1572 -2790
rect -652 -3710 -628 -2790
rect -1596 -3734 -628 -3710
rect -308 -2811 12 -2769
rect -308 -3689 -266 -2811
rect -30 -3689 12 -2811
rect -308 -3731 12 -3689
rect 126 -2790 1094 -2766
rect 126 -3710 150 -2790
rect 1070 -3710 1094 -2790
rect 126 -3734 1094 -3710
rect 1414 -2811 1734 -2769
rect 1414 -3689 1456 -2811
rect 1692 -3689 1734 -2811
rect 1414 -3731 1734 -3689
rect 1848 -2790 2816 -2766
rect 1848 -3710 1872 -2790
rect 2792 -3710 2816 -2790
rect 1848 -3734 2816 -3710
rect 3136 -2811 3456 -2769
rect 3136 -3689 3178 -2811
rect 3414 -3689 3456 -2811
rect 3136 -3731 3456 -3689
rect 3570 -2790 4538 -2766
rect 3570 -3710 3594 -2790
rect 4514 -3710 4538 -2790
rect 3570 -3734 4538 -3710
rect 4858 -2811 5178 -2769
rect 4858 -3689 4900 -2811
rect 5136 -3689 5178 -2811
rect 4858 -3731 5178 -3689
rect -4716 -4066 -4396 -3734
rect -2994 -4066 -2674 -3734
rect -1272 -4066 -952 -3734
rect 450 -4066 770 -3734
rect 2172 -4066 2492 -3734
rect 3894 -4066 4214 -3734
rect -5040 -4090 -4072 -4066
rect -5040 -5010 -5016 -4090
rect -4096 -5010 -4072 -4090
rect -5040 -5034 -4072 -5010
rect -3752 -4111 -3432 -4069
rect -3752 -4989 -3710 -4111
rect -3474 -4989 -3432 -4111
rect -3752 -5031 -3432 -4989
rect -3318 -4090 -2350 -4066
rect -3318 -5010 -3294 -4090
rect -2374 -5010 -2350 -4090
rect -3318 -5034 -2350 -5010
rect -2030 -4111 -1710 -4069
rect -2030 -4989 -1988 -4111
rect -1752 -4989 -1710 -4111
rect -2030 -5031 -1710 -4989
rect -1596 -4090 -628 -4066
rect -1596 -5010 -1572 -4090
rect -652 -5010 -628 -4090
rect -1596 -5034 -628 -5010
rect -308 -4111 12 -4069
rect -308 -4989 -266 -4111
rect -30 -4989 12 -4111
rect -308 -5031 12 -4989
rect 126 -4090 1094 -4066
rect 126 -5010 150 -4090
rect 1070 -5010 1094 -4090
rect 126 -5034 1094 -5010
rect 1414 -4111 1734 -4069
rect 1414 -4989 1456 -4111
rect 1692 -4989 1734 -4111
rect 1414 -5031 1734 -4989
rect 1848 -4090 2816 -4066
rect 1848 -5010 1872 -4090
rect 2792 -5010 2816 -4090
rect 1848 -5034 2816 -5010
rect 3136 -4111 3456 -4069
rect 3136 -4989 3178 -4111
rect 3414 -4989 3456 -4111
rect 3136 -5031 3456 -4989
rect 3570 -4090 4538 -4066
rect 3570 -5010 3594 -4090
rect 4514 -5010 4538 -4090
rect 3570 -5034 4538 -5010
rect 4858 -4111 5178 -4069
rect 4858 -4989 4900 -4111
rect 5136 -4989 5178 -4111
rect 4858 -5031 5178 -4989
rect -4716 -5366 -4396 -5034
rect -2994 -5366 -2674 -5034
rect -1272 -5366 -952 -5034
rect 450 -5366 770 -5034
rect 2172 -5366 2492 -5034
rect 3894 -5366 4214 -5034
rect -5040 -5390 -4072 -5366
rect -5040 -6310 -5016 -5390
rect -4096 -6310 -4072 -5390
rect -5040 -6334 -4072 -6310
rect -3752 -5411 -3432 -5369
rect -3752 -6289 -3710 -5411
rect -3474 -6289 -3432 -5411
rect -3752 -6331 -3432 -6289
rect -3318 -5390 -2350 -5366
rect -3318 -6310 -3294 -5390
rect -2374 -6310 -2350 -5390
rect -3318 -6334 -2350 -6310
rect -2030 -5411 -1710 -5369
rect -2030 -6289 -1988 -5411
rect -1752 -6289 -1710 -5411
rect -2030 -6331 -1710 -6289
rect -1596 -5390 -628 -5366
rect -1596 -6310 -1572 -5390
rect -652 -6310 -628 -5390
rect -1596 -6334 -628 -6310
rect -308 -5411 12 -5369
rect -308 -6289 -266 -5411
rect -30 -6289 12 -5411
rect -308 -6331 12 -6289
rect 126 -5390 1094 -5366
rect 126 -6310 150 -5390
rect 1070 -6310 1094 -5390
rect 126 -6334 1094 -6310
rect 1414 -5411 1734 -5369
rect 1414 -6289 1456 -5411
rect 1692 -6289 1734 -5411
rect 1414 -6331 1734 -6289
rect 1848 -5390 2816 -5366
rect 1848 -6310 1872 -5390
rect 2792 -6310 2816 -5390
rect 1848 -6334 2816 -6310
rect 3136 -5411 3456 -5369
rect 3136 -6289 3178 -5411
rect 3414 -6289 3456 -5411
rect 3136 -6331 3456 -6289
rect 3570 -5390 4538 -5366
rect 3570 -6310 3594 -5390
rect 4514 -6310 4538 -5390
rect 3570 -6334 4538 -6310
rect 4858 -5411 5178 -5369
rect 4858 -6289 4900 -5411
rect 5136 -6289 5178 -5411
rect 4858 -6331 5178 -6289
rect -4716 -6500 -4396 -6334
rect -2994 -6500 -2674 -6334
rect -1272 -6500 -952 -6334
rect 450 -6500 770 -6334
rect 2172 -6500 2492 -6334
rect 3894 -6500 4214 -6334
<< properties >>
string FIXED_BBOX 3454 5250 4654 6450
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 6 ny 10 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 1 ccov 100
<< end >>
