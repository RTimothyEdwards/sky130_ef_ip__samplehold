magic
tech sky130A
magscale 1 2
timestamp 1718242347
<< nwell >>
rect -387 -762 387 762
<< mvpmos >>
rect -129 -464 -29 536
rect 29 -464 129 536
<< mvpdiff >>
rect -187 524 -129 536
rect -187 -452 -175 524
rect -141 -452 -129 524
rect -187 -464 -129 -452
rect -29 524 29 536
rect -29 -452 -17 524
rect 17 -452 29 524
rect -29 -464 29 -452
rect 129 524 187 536
rect 129 -452 141 524
rect 175 -452 187 524
rect 129 -464 187 -452
<< mvpdiffc >>
rect -175 -452 -141 524
rect -17 -452 17 524
rect 141 -452 175 524
<< mvnsubdiff >>
rect -321 684 321 696
rect -321 650 -213 684
rect 213 650 321 684
rect -321 638 321 650
rect -321 588 -263 638
rect -321 -588 -309 588
rect -275 -588 -263 588
rect 263 588 321 638
rect -321 -638 -263 -588
rect 263 -588 275 588
rect 309 -588 321 588
rect 263 -638 321 -588
rect -321 -650 321 -638
rect -321 -684 -213 -650
rect 213 -684 321 -650
rect -321 -696 321 -684
<< mvnsubdiffcont >>
rect -213 650 213 684
rect -309 -588 -275 588
rect 275 -588 309 588
rect -213 -684 213 -650
<< poly >>
rect -129 536 -29 562
rect 29 536 129 562
rect -129 -511 -29 -464
rect -129 -545 -113 -511
rect -45 -545 -29 -511
rect -129 -561 -29 -545
rect 29 -511 129 -464
rect 29 -545 45 -511
rect 113 -545 129 -511
rect 29 -561 129 -545
<< polycont >>
rect -113 -545 -45 -511
rect 45 -545 113 -511
<< locali >>
rect -309 650 -213 684
rect 213 650 309 684
rect -309 588 -275 650
rect 275 588 309 650
rect -175 524 -141 540
rect -175 -468 -141 -452
rect -17 524 17 540
rect -17 -468 17 -452
rect 141 524 175 540
rect 141 -468 175 -452
rect -129 -545 -113 -511
rect -45 -545 -29 -511
rect 29 -545 45 -511
rect 113 -545 129 -511
rect -309 -650 -275 -588
rect 275 -650 309 -588
rect -309 -684 -213 -650
rect 213 -684 309 -650
<< viali >>
rect -175 -452 -141 524
rect -17 -452 17 524
rect 141 -452 175 524
rect -113 -545 -45 -511
rect 45 -545 113 -511
<< metal1 >>
rect -181 524 -135 536
rect -181 -452 -175 524
rect -141 -452 -135 524
rect -181 -464 -135 -452
rect -23 524 23 536
rect -23 -452 -17 524
rect 17 -452 23 524
rect -23 -464 23 -452
rect 135 524 181 536
rect 135 -452 141 524
rect 175 -452 181 524
rect 135 -464 181 -452
rect -125 -511 -33 -505
rect -125 -545 -113 -511
rect -45 -545 -33 -511
rect -125 -551 -33 -545
rect 33 -511 125 -505
rect 33 -545 45 -511
rect 113 -545 125 -511
rect 33 -551 125 -545
<< properties >>
string FIXED_BBOX -292 -667 292 667
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
