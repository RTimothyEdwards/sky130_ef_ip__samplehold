magic
tech sky130A
timestamp 1651947168
<< end >>
