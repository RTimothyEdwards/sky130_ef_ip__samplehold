magic
tech sky130A
magscale 1 2
timestamp 1718242007
<< nwell >>
rect -387 -512 387 512
<< mvpmos >>
rect -129 -214 -29 286
rect 29 -214 129 286
<< mvpdiff >>
rect -187 274 -129 286
rect -187 -202 -175 274
rect -141 -202 -129 274
rect -187 -214 -129 -202
rect -29 274 29 286
rect -29 -202 -17 274
rect 17 -202 29 274
rect -29 -214 29 -202
rect 129 274 187 286
rect 129 -202 141 274
rect 175 -202 187 274
rect 129 -214 187 -202
<< mvpdiffc >>
rect -175 -202 -141 274
rect -17 -202 17 274
rect 141 -202 175 274
<< mvnsubdiff >>
rect -321 434 321 446
rect -321 400 -213 434
rect 213 400 321 434
rect -321 388 321 400
rect -321 338 -263 388
rect -321 -338 -309 338
rect -275 -338 -263 338
rect 263 338 321 388
rect -321 -388 -263 -338
rect 263 -338 275 338
rect 309 -338 321 338
rect 263 -388 321 -338
rect -321 -400 321 -388
rect -321 -434 -213 -400
rect 213 -434 321 -400
rect -321 -446 321 -434
<< mvnsubdiffcont >>
rect -213 400 213 434
rect -309 -338 -275 338
rect 275 -338 309 338
rect -213 -434 213 -400
<< poly >>
rect -129 286 -29 312
rect 29 286 129 312
rect -129 -261 -29 -214
rect -129 -295 -113 -261
rect -45 -295 -29 -261
rect -129 -311 -29 -295
rect 29 -261 129 -214
rect 29 -295 45 -261
rect 113 -295 129 -261
rect 29 -311 129 -295
<< polycont >>
rect -113 -295 -45 -261
rect 45 -295 113 -261
<< locali >>
rect -309 400 -213 434
rect 213 400 309 434
rect -309 338 -275 400
rect 275 338 309 400
rect -175 274 -141 290
rect -175 -218 -141 -202
rect -17 274 17 290
rect -17 -218 17 -202
rect 141 274 175 290
rect 141 -218 175 -202
rect -129 -295 -113 -261
rect -45 -295 -29 -261
rect 29 -295 45 -261
rect 113 -295 129 -261
rect -309 -400 -275 -338
rect 275 -400 309 -338
rect -309 -434 -213 -400
rect 213 -434 309 -400
<< viali >>
rect -175 -202 -141 274
rect -17 -202 17 274
rect 141 -202 175 274
rect -113 -295 -45 -261
rect 45 -295 113 -261
<< metal1 >>
rect -181 274 -135 286
rect -181 -202 -175 274
rect -141 -202 -135 274
rect -181 -214 -135 -202
rect -23 274 23 286
rect -23 -202 -17 274
rect 17 -202 23 274
rect -23 -214 23 -202
rect 135 274 181 286
rect 135 -202 141 274
rect 175 -202 181 274
rect 135 -214 181 -202
rect -125 -261 -33 -255
rect -125 -295 -113 -261
rect -45 -295 -33 -261
rect -125 -301 -33 -295
rect 33 -261 125 -255
rect 33 -295 45 -261
rect 113 -295 125 -261
rect 33 -301 125 -295
<< properties >>
string FIXED_BBOX -292 -417 292 417
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2.5 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
