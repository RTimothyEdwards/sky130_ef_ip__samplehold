magic
tech sky130A
magscale 1 2
timestamp 1652200182
<< dnwell >>
rect 410 -2200 2434 1630
<< nwell >>
rect 301 1424 2543 1830
rect 301 482 616 1424
rect 2228 482 2543 1424
rect 301 373 2543 482
rect 301 -1994 616 373
rect 1957 -297 2543 373
rect 2228 -1994 2543 -297
rect 301 -2311 2543 -1994
<< mvnsubdiff >>
rect 367 1744 2477 1764
rect 367 1710 447 1744
rect 2397 1710 2477 1744
rect 367 1690 2477 1710
rect 367 1684 441 1690
rect 367 -2163 387 1684
rect 421 -2163 441 1684
rect 367 -2169 441 -2163
rect 2403 1684 2477 1690
rect 2403 -2163 2423 1684
rect 2457 -2163 2477 1684
rect 2403 -2169 2477 -2163
rect 367 -2189 2477 -2169
rect 367 -2223 447 -2189
rect 2397 -2223 2477 -2189
rect 367 -2243 2477 -2223
<< mvnsubdiffcont >>
rect 447 1710 2397 1744
rect 387 -2163 421 1684
rect 2423 -2163 2457 1684
rect 447 -2223 2397 -2189
<< locali >>
rect 387 1710 447 1744
rect 2397 1710 2457 1744
rect 387 1684 2457 1710
rect 421 1621 2423 1684
rect 421 482 571 1621
rect 616 556 768 1376
rect 1169 1355 1343 1377
rect 1169 674 1221 1355
rect 1297 674 1343 1355
rect 1169 556 1343 674
rect 1753 1357 2255 1377
rect 1753 676 1802 1357
rect 1878 847 2255 1357
rect 1878 676 1927 847
rect 1753 556 1927 676
rect 2164 556 2255 847
rect 2325 482 2423 1621
rect 421 342 2423 482
rect 421 -158 712 342
rect 1870 -158 2423 342
rect 421 -185 2423 -158
rect 421 -358 537 -185
rect 2337 -358 2423 -185
rect 421 -374 2423 -358
rect 421 -894 712 -374
rect 2140 -894 2423 -374
rect 421 -988 2423 -894
rect 421 -1828 528 -988
rect 599 -1155 2235 -1066
rect 599 -1870 714 -1155
rect 2120 -1870 2235 -1155
rect 2302 -1821 2423 -988
rect 471 -1911 2378 -1870
rect 471 -2081 582 -1911
rect 2327 -2081 2378 -1911
rect 471 -2143 2378 -2081
rect 387 -2189 421 -2163
rect 2423 -2189 2457 -2163
rect 387 -2223 447 -2189
rect 2397 -2223 2457 -2189
<< viali >>
rect 1221 674 1297 1355
rect 1802 676 1878 1357
rect 537 -358 2337 -185
rect 582 -2081 2327 -1911
<< metal1 >>
rect 393 1541 2463 1563
rect 393 1322 544 1541
rect 842 1357 2463 1541
rect 842 1355 1802 1357
rect 842 1322 1221 1355
rect 393 1306 1221 1322
rect 824 764 888 1306
rect 340 619 540 690
rect 943 619 980 1231
rect 340 567 894 619
rect 972 567 980 619
rect 340 490 540 567
rect 943 401 980 567
rect 1052 502 1101 1172
rect 1211 674 1221 1306
rect 1297 1306 1802 1355
rect 1297 674 1308 1306
rect 1406 760 1470 1306
rect 1211 659 1308 674
rect 1534 502 1571 1232
rect 1052 453 1571 502
rect 909 364 1099 401
rect 909 200 946 364
rect 1062 200 1099 364
rect 793 138 866 153
rect 793 -46 803 138
rect 857 -46 866 138
rect 793 -59 866 -46
rect 964 -92 1036 156
rect 1158 139 1207 453
rect 1534 401 1571 453
rect 1620 500 1669 1171
rect 1791 676 1802 1306
rect 1878 1306 2463 1357
rect 1878 676 1888 1306
rect 1791 664 1888 676
rect 2009 619 2080 739
rect 2009 561 2080 567
rect 1620 451 1792 500
rect 1490 364 1680 401
rect 1490 200 1527 364
rect 1643 200 1680 364
rect 1201 -45 1207 139
rect 1158 -57 1207 -45
rect 1375 140 1448 151
rect 1375 -44 1382 140
rect 1436 -44 1448 140
rect 1375 -61 1448 -44
rect 1552 -92 1624 151
rect 1743 140 1792 451
rect 1786 -44 1792 140
rect 1743 -59 1792 -44
rect 326 -185 2478 -92
rect 326 -358 537 -185
rect 2337 -358 2478 -185
rect 326 -368 2478 -358
rect 904 -449 959 -397
rect 1040 -449 1046 -397
rect 904 -453 1046 -449
rect 745 -642 867 -636
rect 745 -695 751 -642
rect 860 -695 867 -642
rect 745 -701 867 -695
rect 904 -867 939 -453
rect 1370 -455 1376 -402
rect 1457 -455 1525 -402
rect 1370 -458 1525 -455
rect 1190 -501 1292 -495
rect 1190 -585 1196 -501
rect 1286 -585 1292 -501
rect 1190 -591 1292 -585
rect 977 -641 1099 -635
rect 977 -694 984 -641
rect 1093 -694 1099 -641
rect 977 -700 1099 -694
rect 1350 -714 1356 -648
rect 1446 -714 1452 -648
rect 1489 -749 1525 -458
rect 1562 -501 1664 -495
rect 1562 -585 1568 -501
rect 1658 -585 1664 -501
rect 1755 -511 1876 -505
rect 1755 -564 1761 -511
rect 1870 -564 1876 -511
rect 1755 -570 1876 -564
rect 1988 -511 2109 -505
rect 1988 -564 1994 -511
rect 2103 -564 2109 -511
rect 1988 -570 2109 -564
rect 1562 -591 1664 -585
rect 1334 -779 1685 -749
rect 1334 -785 1623 -779
rect 1617 -839 1623 -785
rect 1679 -839 1685 -779
rect 1913 -867 1948 -760
rect 904 -915 1948 -867
rect 2209 -776 2526 -576
rect 2209 -782 2393 -776
rect 314 -968 891 -964
rect 314 -1160 735 -968
rect 885 -1160 891 -968
rect 314 -1164 891 -1160
rect 1051 -1045 1128 -1037
rect 1051 -1107 1128 -1101
rect 1051 -1261 1087 -1107
rect 894 -1289 1087 -1261
rect 1479 -1264 1515 -915
rect 1728 -1045 1805 -1039
rect 1728 -1109 1805 -1101
rect 887 -1297 1087 -1289
rect 740 -1348 856 -1342
rect 740 -1485 746 -1348
rect 850 -1485 856 -1348
rect 740 -1491 856 -1485
rect 887 -1784 923 -1297
rect 1322 -1300 1515 -1264
rect 1756 -1262 1792 -1109
rect 2209 -1226 2217 -782
rect 2387 -1226 2393 -782
rect 2209 -1236 2393 -1226
rect 1756 -1298 1949 -1262
rect 967 -1348 1083 -1342
rect 967 -1485 973 -1348
rect 1077 -1485 1083 -1348
rect 967 -1491 1083 -1485
rect 1323 -1358 1440 -1352
rect 1323 -1482 1329 -1358
rect 1434 -1482 1440 -1358
rect 1323 -1488 1440 -1482
rect 1166 -1587 1282 -1581
rect 1166 -1724 1172 -1587
rect 1276 -1724 1282 -1587
rect 1166 -1730 1282 -1724
rect 1479 -1773 1515 -1300
rect 1552 -1587 1668 -1581
rect 1552 -1724 1558 -1587
rect 1662 -1724 1668 -1587
rect 1552 -1730 1668 -1724
rect 1750 -1587 1866 -1581
rect 1750 -1724 1756 -1587
rect 1860 -1724 1866 -1587
rect 1750 -1730 1866 -1724
rect 1347 -1809 1515 -1773
rect 1910 -1786 1946 -1298
rect 1978 -1587 2094 -1581
rect 1978 -1724 1984 -1587
rect 2088 -1724 2094 -1587
rect 1978 -1730 2094 -1724
rect 328 -1879 2515 -1870
rect 328 -2098 542 -1879
rect 840 -1911 2515 -1879
rect 2327 -2081 2515 -1911
rect 840 -2098 2515 -2081
rect 328 -2105 2515 -2098
<< via1 >>
rect 544 1322 842 1541
rect 894 567 972 619
rect 803 -46 857 138
rect 2009 567 2080 619
rect 1147 -45 1201 139
rect 1382 -44 1436 140
rect 1732 -44 1786 140
rect 959 -449 1040 -397
rect 751 -695 860 -642
rect 1376 -455 1457 -402
rect 1196 -585 1286 -501
rect 984 -694 1093 -641
rect 1356 -714 1446 -648
rect 1568 -585 1658 -501
rect 1761 -564 1870 -511
rect 1994 -564 2103 -511
rect 1623 -839 1679 -779
rect 735 -1160 885 -968
rect 1051 -1101 1128 -1045
rect 1728 -1101 1805 -1045
rect 746 -1485 850 -1348
rect 2217 -1226 2387 -782
rect 973 -1485 1077 -1348
rect 1329 -1482 1434 -1358
rect 1172 -1724 1276 -1587
rect 1558 -1724 1662 -1587
rect 1756 -1724 1860 -1587
rect 1984 -1724 2088 -1587
rect 542 -1911 840 -1879
rect 542 -2081 582 -1911
rect 582 -2081 840 -1911
rect 542 -2098 840 -2081
<< metal2 >>
rect 529 1541 867 1556
rect 529 1322 544 1541
rect 842 1322 867 1541
rect 529 1306 867 1322
rect 529 -1870 660 1306
rect 886 567 894 619
rect 972 567 2009 619
rect 2080 567 2087 619
rect 795 139 1207 141
rect 795 138 1147 139
rect 795 -46 803 138
rect 857 -45 1147 138
rect 1201 -45 1207 139
rect 857 -46 1207 -45
rect 795 -47 1207 -46
rect 1376 140 1792 142
rect 1376 -44 1382 140
rect 1436 -44 1732 140
rect 1786 -44 1792 140
rect 1376 -46 1792 -44
rect 959 -397 1040 -47
rect 959 -455 1040 -449
rect 1376 -402 1457 -46
rect 1376 -461 1457 -455
rect 736 -501 2393 -489
rect 736 -585 1196 -501
rect 1286 -585 1568 -501
rect 1658 -511 2393 -501
rect 1658 -564 1761 -511
rect 1870 -564 1994 -511
rect 2103 -564 2393 -511
rect 1658 -585 2393 -564
rect 736 -593 2393 -585
rect 732 -641 2127 -634
rect 732 -642 984 -641
rect 732 -695 751 -642
rect 860 -694 984 -642
rect 1093 -648 2127 -641
rect 1093 -694 1356 -648
rect 860 -695 1356 -694
rect 732 -714 1356 -695
rect 1446 -714 2127 -648
rect 732 -738 2127 -714
rect 732 -968 891 -738
rect 732 -1160 735 -968
rect 885 -1160 891 -968
rect 1623 -779 1679 -772
rect 1623 -1045 1679 -839
rect 2209 -782 2393 -593
rect 1043 -1101 1051 -1045
rect 1128 -1101 1728 -1045
rect 1805 -1101 1816 -1045
rect 732 -1313 891 -1160
rect 2209 -1226 2217 -782
rect 2387 -1226 2393 -782
rect 732 -1348 2122 -1313
rect 732 -1485 746 -1348
rect 850 -1485 973 -1348
rect 1077 -1358 2122 -1348
rect 1077 -1482 1329 -1358
rect 1434 -1482 2122 -1358
rect 1077 -1485 2122 -1482
rect 732 -1497 2122 -1485
rect 2209 -1558 2393 -1226
rect 733 -1587 2393 -1558
rect 733 -1724 1172 -1587
rect 1276 -1724 1558 -1587
rect 1662 -1724 1756 -1587
rect 1860 -1724 1984 -1587
rect 2088 -1724 2393 -1587
rect 733 -1742 2393 -1724
rect 529 -1879 849 -1870
rect 529 -2098 542 -1879
rect 840 -2098 849 -1879
rect 529 -2105 849 -2098
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XD1 paramcells
timestamp 1652200182
transform 1 0 2045 0 -1 703
box -183 -183 183 183
use sky130_fd_pr__nfet_g5v0d10v5_EJGQFX  XM1 paramcells
timestamp 1652200182
transform -1 0 1417 0 1 -1536
box -357 -458 357 458
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM3 paramcells
timestamp 1652200182
transform -1 0 907 0 1 -1536
box -278 -458 278 458
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM4 paramcells
timestamp 1652200182
transform 1 0 1427 0 1 -638
box -387 -362 387 362
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM5
timestamp 1652200182
transform 1 0 1927 0 1 -1536
box -278 -458 278 458
use sky130_fd_pr__pfet_g5v0d10v5_U6NWY6  XM6 paramcells
timestamp 1652200182
transform 1 0 1932 0 1 -638
box -308 -362 308 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM7
timestamp 1652200182
transform 1 0 1001 0 -1 82
box -387 -362 387 362
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM8
timestamp 1652200182
transform 1 0 964 0 -1 966
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM10
timestamp 1652200182
transform 1 0 1546 0 -1 966
box -278 -458 278 458
use sky130_fd_pr__pfet_g5v0d10v5_U6NWY6  sky130_fd_pr__pfet_g5v0d10v5_U6NWY6_0
timestamp 1652200182
transform 1 0 922 0 1 -638
box -308 -362 308 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  sky130_fd_pr__pfet_g5v0d10v5_U62SY6_0
timestamp 1652200182
transform 1 0 1585 0 -1 82
box -387 -362 387 362
<< labels >>
flabel metal1 314 -1164 514 -964 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal1 2326 -776 2526 -576 0 FreeSans 256 0 0 0 out
port 3 nsew
flabel metal1 326 -352 526 -152 0 FreeSans 256 0 0 0 vdd
port 5 nsew
flabel metal1 336 -2091 536 -1891 0 FreeSans 256 0 0 0 vss
port 2 nsew
flabel metal1 340 490 540 690 0 FreeSans 256 0 0 0 hold
port 1 nsew
flabel metal1 1271 478 1271 478 0 FreeSans 320 0 0 0 holdb
flabel metal1 1705 473 1705 473 0 FreeSans 320 0 0 0 holdp
<< end >>
