magic
tech sky130A
magscale 1 2
timestamp 1651944383
<< error_p >>
rect -1792 2431 -1732 2550
rect -1712 2431 -1652 2550
rect -1916 1469 -1652 2431
rect -1792 1350 -1732 1469
rect -1712 1350 -1652 1469
rect -1596 1466 -1390 2434
rect -70 2431 -10 2550
rect 10 2431 70 2550
rect -194 1469 70 2431
rect -70 1350 -10 1469
rect 10 1350 70 1469
rect 126 1466 332 2434
rect 1652 2431 1712 2550
rect 1732 2431 1792 2550
rect 1528 1469 1792 2431
rect 1652 1350 1712 1469
rect 1732 1350 1792 1469
rect 1848 1466 2054 2434
rect -1792 1131 -1732 1250
rect -1712 1131 -1652 1250
rect -1916 169 -1652 1131
rect -1792 50 -1732 169
rect -1712 50 -1652 169
rect -1596 166 -1390 1134
rect -70 1131 -10 1250
rect 10 1131 70 1250
rect -194 169 70 1131
rect -70 50 -10 169
rect 10 50 70 169
rect 126 166 332 1134
rect 1652 1131 1712 1250
rect 1732 1131 1792 1250
rect 1528 169 1792 1131
rect 1652 50 1712 169
rect 1732 50 1792 169
rect 1848 166 2054 1134
rect -1792 -169 -1732 -50
rect -1712 -169 -1652 -50
rect -1916 -1131 -1652 -169
rect -1792 -1250 -1732 -1131
rect -1712 -1250 -1652 -1131
rect -1596 -1134 -1390 -166
rect -70 -169 -10 -50
rect 10 -169 70 -50
rect -194 -1131 70 -169
rect -70 -1250 -10 -1131
rect 10 -1250 70 -1131
rect 126 -1134 332 -166
rect 1652 -169 1712 -50
rect 1732 -169 1792 -50
rect 1528 -1131 1792 -169
rect 1652 -1250 1712 -1131
rect 1732 -1250 1792 -1131
rect 1848 -1134 2054 -166
rect -1792 -1469 -1732 -1350
rect -1712 -1469 -1652 -1350
rect -1916 -2431 -1652 -1469
rect -1792 -2550 -1732 -2431
rect -1712 -2550 -1652 -2431
rect -1596 -2434 -1390 -1466
rect -70 -1469 -10 -1350
rect 10 -1469 70 -1350
rect -194 -2431 70 -1469
rect -70 -2550 -10 -2431
rect 10 -2550 70 -2431
rect 126 -2434 332 -1466
rect 1652 -1469 1712 -1350
rect 1732 -1469 1792 -1350
rect 1528 -2431 1792 -1469
rect 1652 -2550 1712 -2431
rect 1732 -2550 1792 -2431
rect 1848 -2434 2054 -1466
<< metal4 >>
rect -3434 2389 -1732 2550
rect -3434 1511 -1988 2389
rect -1752 1511 -1732 2389
rect -3434 1350 -1732 1511
rect -1712 2389 -10 2550
rect -1712 1511 -266 2389
rect -30 1511 -10 2389
rect -1712 1350 -10 1511
rect 10 2389 1712 2550
rect 10 1511 1456 2389
rect 1692 1511 1712 2389
rect 10 1350 1712 1511
rect 1732 2389 3434 2550
rect 1732 1511 3178 2389
rect 3414 1511 3434 2389
rect 1732 1350 3434 1511
rect -3434 1089 -1732 1250
rect -3434 211 -1988 1089
rect -1752 211 -1732 1089
rect -3434 50 -1732 211
rect -1712 1089 -10 1250
rect -1712 211 -266 1089
rect -30 211 -10 1089
rect -1712 50 -10 211
rect 10 1089 1712 1250
rect 10 211 1456 1089
rect 1692 211 1712 1089
rect 10 50 1712 211
rect 1732 1089 3434 1250
rect 1732 211 3178 1089
rect 3414 211 3434 1089
rect 1732 50 3434 211
rect -3434 -211 -1732 -50
rect -3434 -1089 -1988 -211
rect -1752 -1089 -1732 -211
rect -3434 -1250 -1732 -1089
rect -1712 -211 -10 -50
rect -1712 -1089 -266 -211
rect -30 -1089 -10 -211
rect -1712 -1250 -10 -1089
rect 10 -211 1712 -50
rect 10 -1089 1456 -211
rect 1692 -1089 1712 -211
rect 10 -1250 1712 -1089
rect 1732 -211 3434 -50
rect 1732 -1089 3178 -211
rect 3414 -1089 3434 -211
rect 1732 -1250 3434 -1089
rect -3434 -1511 -1732 -1350
rect -3434 -2389 -1988 -1511
rect -1752 -2389 -1732 -1511
rect -3434 -2550 -1732 -2389
rect -1712 -1511 -10 -1350
rect -1712 -2389 -266 -1511
rect -30 -2389 -10 -1511
rect -1712 -2550 -10 -2389
rect 10 -1511 1712 -1350
rect 10 -2389 1456 -1511
rect 1692 -2389 1712 -1511
rect 10 -2550 1712 -2389
rect 1732 -1511 3434 -1350
rect 1732 -2389 3178 -1511
rect 3414 -2389 3434 -1511
rect 1732 -2550 3434 -2389
<< via4 >>
rect -1988 1511 -1752 2389
rect -266 1511 -30 2389
rect 1456 1511 1692 2389
rect 3178 1511 3414 2389
rect -1988 211 -1752 1089
rect -266 211 -30 1089
rect 1456 211 1692 1089
rect 3178 211 3414 1089
rect -1988 -1089 -1752 -211
rect -266 -1089 -30 -211
rect 1456 -1089 1692 -211
rect 3178 -1089 3414 -211
rect -1988 -2389 -1752 -1511
rect -266 -2389 -30 -1511
rect 1456 -2389 1692 -1511
rect 3178 -2389 3414 -1511
<< mimcap2 >>
rect -3334 2410 -2334 2450
rect -3334 1490 -3294 2410
rect -2374 1490 -2334 2410
rect -3334 1450 -2334 1490
rect -1612 2410 -612 2450
rect -1612 1490 -1572 2410
rect -652 1490 -612 2410
rect -1612 1450 -612 1490
rect 110 2410 1110 2450
rect 110 1490 150 2410
rect 1070 1490 1110 2410
rect 110 1450 1110 1490
rect 1832 2410 2832 2450
rect 1832 1490 1872 2410
rect 2792 1490 2832 2410
rect 1832 1450 2832 1490
rect -3334 1110 -2334 1150
rect -3334 190 -3294 1110
rect -2374 190 -2334 1110
rect -3334 150 -2334 190
rect -1612 1110 -612 1150
rect -1612 190 -1572 1110
rect -652 190 -612 1110
rect -1612 150 -612 190
rect 110 1110 1110 1150
rect 110 190 150 1110
rect 1070 190 1110 1110
rect 110 150 1110 190
rect 1832 1110 2832 1150
rect 1832 190 1872 1110
rect 2792 190 2832 1110
rect 1832 150 2832 190
rect -3334 -190 -2334 -150
rect -3334 -1110 -3294 -190
rect -2374 -1110 -2334 -190
rect -3334 -1150 -2334 -1110
rect -1612 -190 -612 -150
rect -1612 -1110 -1572 -190
rect -652 -1110 -612 -190
rect -1612 -1150 -612 -1110
rect 110 -190 1110 -150
rect 110 -1110 150 -190
rect 1070 -1110 1110 -190
rect 110 -1150 1110 -1110
rect 1832 -190 2832 -150
rect 1832 -1110 1872 -190
rect 2792 -1110 2832 -190
rect 1832 -1150 2832 -1110
rect -3334 -1490 -2334 -1450
rect -3334 -2410 -3294 -1490
rect -2374 -2410 -2334 -1490
rect -3334 -2450 -2334 -2410
rect -1612 -1490 -612 -1450
rect -1612 -2410 -1572 -1490
rect -652 -2410 -612 -1490
rect -1612 -2450 -612 -2410
rect 110 -1490 1110 -1450
rect 110 -2410 150 -1490
rect 1070 -2410 1110 -1490
rect 110 -2450 1110 -2410
rect 1832 -1490 2832 -1450
rect 1832 -2410 1872 -1490
rect 2792 -2410 2832 -1490
rect 1832 -2450 2832 -2410
<< mimcap2contact >>
rect -3294 1490 -2374 2410
rect -1572 1490 -652 2410
rect 150 1490 1070 2410
rect 1872 1490 2792 2410
rect -3294 190 -2374 1110
rect -1572 190 -652 1110
rect 150 190 1070 1110
rect 1872 190 2792 1110
rect -3294 -1110 -2374 -190
rect -1572 -1110 -652 -190
rect 150 -1110 1070 -190
rect 1872 -1110 2792 -190
rect -3294 -2410 -2374 -1490
rect -1572 -2410 -652 -1490
rect 150 -2410 1070 -1490
rect 1872 -2410 2792 -1490
<< metal5 >>
rect -2994 2434 -2674 2600
rect -1272 2434 -952 2600
rect 450 2434 770 2600
rect 2172 2434 2492 2600
rect -3318 2410 -2350 2434
rect -3318 1490 -3294 2410
rect -2374 1490 -2350 2410
rect -3318 1466 -2350 1490
rect -2030 2389 -1710 2431
rect -2030 1511 -1988 2389
rect -1752 1511 -1710 2389
rect -2030 1469 -1710 1511
rect -1596 2410 -628 2434
rect -1596 1490 -1572 2410
rect -652 1490 -628 2410
rect -1596 1466 -628 1490
rect -308 2389 12 2431
rect -308 1511 -266 2389
rect -30 1511 12 2389
rect -308 1469 12 1511
rect 126 2410 1094 2434
rect 126 1490 150 2410
rect 1070 1490 1094 2410
rect 126 1466 1094 1490
rect 1414 2389 1734 2431
rect 1414 1511 1456 2389
rect 1692 1511 1734 2389
rect 1414 1469 1734 1511
rect 1848 2410 2816 2434
rect 1848 1490 1872 2410
rect 2792 1490 2816 2410
rect 1848 1466 2816 1490
rect 3136 2389 3456 2431
rect 3136 1511 3178 2389
rect 3414 1511 3456 2389
rect 3136 1469 3456 1511
rect -2994 1134 -2674 1466
rect -1272 1134 -952 1466
rect 450 1134 770 1466
rect 2172 1134 2492 1466
rect -3318 1110 -2350 1134
rect -3318 190 -3294 1110
rect -2374 190 -2350 1110
rect -3318 166 -2350 190
rect -2030 1089 -1710 1131
rect -2030 211 -1988 1089
rect -1752 211 -1710 1089
rect -2030 169 -1710 211
rect -1596 1110 -628 1134
rect -1596 190 -1572 1110
rect -652 190 -628 1110
rect -1596 166 -628 190
rect -308 1089 12 1131
rect -308 211 -266 1089
rect -30 211 12 1089
rect -308 169 12 211
rect 126 1110 1094 1134
rect 126 190 150 1110
rect 1070 190 1094 1110
rect 126 166 1094 190
rect 1414 1089 1734 1131
rect 1414 211 1456 1089
rect 1692 211 1734 1089
rect 1414 169 1734 211
rect 1848 1110 2816 1134
rect 1848 190 1872 1110
rect 2792 190 2816 1110
rect 1848 166 2816 190
rect 3136 1089 3456 1131
rect 3136 211 3178 1089
rect 3414 211 3456 1089
rect 3136 169 3456 211
rect -2994 -166 -2674 166
rect -1272 -166 -952 166
rect 450 -166 770 166
rect 2172 -166 2492 166
rect -3318 -190 -2350 -166
rect -3318 -1110 -3294 -190
rect -2374 -1110 -2350 -190
rect -3318 -1134 -2350 -1110
rect -2030 -211 -1710 -169
rect -2030 -1089 -1988 -211
rect -1752 -1089 -1710 -211
rect -2030 -1131 -1710 -1089
rect -1596 -190 -628 -166
rect -1596 -1110 -1572 -190
rect -652 -1110 -628 -190
rect -1596 -1134 -628 -1110
rect -308 -211 12 -169
rect -308 -1089 -266 -211
rect -30 -1089 12 -211
rect -308 -1131 12 -1089
rect 126 -190 1094 -166
rect 126 -1110 150 -190
rect 1070 -1110 1094 -190
rect 126 -1134 1094 -1110
rect 1414 -211 1734 -169
rect 1414 -1089 1456 -211
rect 1692 -1089 1734 -211
rect 1414 -1131 1734 -1089
rect 1848 -190 2816 -166
rect 1848 -1110 1872 -190
rect 2792 -1110 2816 -190
rect 1848 -1134 2816 -1110
rect 3136 -211 3456 -169
rect 3136 -1089 3178 -211
rect 3414 -1089 3456 -211
rect 3136 -1131 3456 -1089
rect -2994 -1466 -2674 -1134
rect -1272 -1466 -952 -1134
rect 450 -1466 770 -1134
rect 2172 -1466 2492 -1134
rect -3318 -1490 -2350 -1466
rect -3318 -2410 -3294 -1490
rect -2374 -2410 -2350 -1490
rect -3318 -2434 -2350 -2410
rect -2030 -1511 -1710 -1469
rect -2030 -2389 -1988 -1511
rect -1752 -2389 -1710 -1511
rect -2030 -2431 -1710 -2389
rect -1596 -1490 -628 -1466
rect -1596 -2410 -1572 -1490
rect -652 -2410 -628 -1490
rect -1596 -2434 -628 -2410
rect -308 -1511 12 -1469
rect -308 -2389 -266 -1511
rect -30 -2389 12 -1511
rect -308 -2431 12 -2389
rect 126 -1490 1094 -1466
rect 126 -2410 150 -1490
rect 1070 -2410 1094 -1490
rect 126 -2434 1094 -2410
rect 1414 -1511 1734 -1469
rect 1414 -2389 1456 -1511
rect 1692 -2389 1734 -1511
rect 1414 -2431 1734 -2389
rect 1848 -1490 2816 -1466
rect 1848 -2410 1872 -1490
rect 2792 -2410 2816 -1490
rect 1848 -2434 2816 -2410
rect 3136 -1511 3456 -1469
rect 3136 -2389 3178 -1511
rect 3414 -2389 3456 -1511
rect 3136 -2431 3456 -2389
rect -2994 -2600 -2674 -2434
rect -1272 -2600 -952 -2434
rect 450 -2600 770 -2434
rect 2172 -2600 2492 -2434
<< properties >>
string FIXED_BBOX 1732 1350 2932 2550
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 1 ccov 100
<< end >>
