magic
tech sky130A
magscale 1 2
timestamp 1651944383
<< error_p >>
rect -296 273 -263 385
rect -168 333 -141 353
rect -129 333 -29 391
rect -17 333 17 353
rect 29 333 129 391
rect 141 333 168 353
rect -187 331 -175 333
rect -168 331 168 333
rect 175 331 187 333
rect -242 306 -187 331
rect -175 327 -141 331
rect -129 327 -104 331
rect -54 327 -29 331
rect -17 327 17 331
rect 29 327 54 331
rect 104 327 129 331
rect 141 327 175 331
rect -242 285 -209 306
rect -242 273 -196 285
rect -183 273 183 327
rect 187 306 242 331
rect 209 285 242 306
rect 196 273 242 285
rect 263 273 296 385
rect -324 -273 -321 273
rect -296 -273 -196 273
rect -175 -251 -162 273
rect -129 213 -29 273
rect -129 -213 -124 213
rect -30 197 -29 198
rect -17 197 17 228
rect 29 213 129 273
rect 29 197 30 198
rect 34 197 81 213
rect -29 191 81 197
rect -44 147 81 191
rect -44 137 -17 147
rect 17 137 44 147
rect -18 100 -17 101
rect 17 100 43 137
rect -17 99 -16 100
rect 16 99 17 100
rect -107 88 -51 99
rect 51 88 107 99
rect -96 -88 -51 88
rect 62 -88 107 88
rect -17 -100 -16 -99
rect 16 -100 17 -99
rect -18 -101 -17 -100
rect -44 -147 -17 -137
rect 17 -147 81 -100
rect -44 -181 81 -147
rect -44 -191 44 -181
rect -29 -197 43 -191
rect -30 -198 -29 -197
rect 29 -198 30 -197
rect 124 -213 129 213
rect -175 -271 -141 -251
rect -129 -271 -29 -213
rect -17 -271 17 -251
rect 29 -271 129 -213
rect 162 -251 175 273
rect 141 -271 175 -251
rect -184 -273 184 -271
rect 196 -273 296 273
rect 321 -273 324 273
rect -296 -385 -263 -273
rect -242 -285 -196 -273
rect -175 -277 -141 -273
rect -129 -277 -104 -273
rect -54 -277 -29 -273
rect -17 -277 17 -273
rect 29 -277 54 -273
rect 104 -277 129 -273
rect 141 -277 175 -273
rect -242 -306 -209 -285
rect -242 -331 -187 -306
rect -183 -331 183 -277
rect 196 -285 242 -273
rect 209 -306 242 -285
rect 187 -331 242 -306
rect -129 -391 -29 -331
rect 29 -391 129 -331
rect 263 -385 296 -273
<< nwell >>
rect -387 -797 387 797
<< mvpmos >>
rect -129 331 -29 500
rect 29 331 129 500
rect -129 197 -29 273
rect 29 197 129 273
rect -129 181 -17 197
rect 17 181 129 197
rect -129 147 -34 181
rect 34 147 129 181
rect -129 100 -17 147
rect 17 100 129 147
rect -129 88 129 100
rect -129 -88 -96 88
rect -62 -88 62 88
rect 96 -88 129 88
rect -129 -100 129 -88
rect -129 -147 -17 -100
rect 17 -147 129 -100
rect -129 -181 -34 -147
rect 34 -181 129 -147
rect -129 -197 -17 -181
rect 17 -197 129 -181
rect -129 -273 -29 -197
rect 29 -273 129 -197
rect -129 -500 -29 -331
rect 29 -500 129 -331
<< mvpdiff >>
rect -187 488 -129 500
rect -187 331 -175 488
rect -141 331 -129 488
rect -29 488 29 500
rect -29 331 -17 488
rect 17 331 29 488
rect 129 488 187 500
rect 129 331 141 488
rect 175 331 187 488
rect -184 -273 -175 273
rect -141 -273 -129 273
rect -29 197 -17 273
rect 17 197 29 273
rect -29 -273 -17 -197
rect 17 -273 29 -197
rect 129 -273 141 273
rect 175 -273 184 273
rect -187 -488 -175 -331
rect -141 -488 -129 -331
rect -187 -500 -129 -488
rect -29 -488 -17 -331
rect 17 -488 29 -331
rect -29 -500 29 -488
rect 129 -488 141 -331
rect 175 -488 187 -331
rect 129 -500 187 -488
<< mvpdiffc >>
rect -175 331 -141 488
rect -17 331 17 488
rect 141 331 175 488
rect -175 -273 -141 273
rect -17 197 17 273
rect -96 -88 -62 88
rect 62 -88 96 88
rect -17 -273 17 -197
rect 141 -273 175 273
rect -175 -488 -141 -331
rect -17 -488 17 -331
rect 141 -488 175 -331
<< mvnsubdiff >>
rect -321 719 321 731
rect -321 685 -213 719
rect 213 685 321 719
rect -321 673 321 685
rect -321 623 -263 673
rect -321 -623 -309 623
rect -275 -623 -263 623
rect 263 623 321 673
rect -242 319 242 331
rect -242 285 -134 319
rect 134 285 242 319
rect -242 273 242 285
rect -242 223 -184 273
rect -242 -223 -230 223
rect -196 -223 -184 223
rect -242 -273 -184 -223
rect 184 223 242 273
rect 184 -223 196 223
rect 230 -223 242 223
rect 184 -273 242 -223
rect -242 -285 242 -273
rect -242 -319 -134 -285
rect 134 -319 242 -285
rect -242 -331 242 -319
rect -321 -673 -263 -623
rect 263 -623 275 623
rect 309 -623 321 623
rect 263 -673 321 -623
rect -321 -685 321 -673
rect -321 -719 -213 -685
rect 213 -719 321 -685
rect -321 -731 321 -719
<< mvnsubdiffcont >>
rect -213 685 213 719
rect -309 -623 -275 623
rect -134 285 134 319
rect -230 -223 -196 223
rect 196 -223 230 223
rect -134 -319 134 -285
rect 275 -623 309 623
rect -213 -719 213 -685
<< poly >>
rect -129 581 -29 597
rect -129 547 -113 581
rect -45 547 -29 581
rect -129 500 -29 547
rect 29 581 129 597
rect 29 547 45 581
rect 113 547 129 581
rect 29 500 129 547
rect -17 181 17 197
rect -17 100 17 147
rect -17 -147 17 -100
rect -17 -197 17 -181
rect -129 -547 -29 -500
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect -129 -597 -29 -581
rect 29 -547 129 -500
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 29 -597 129 -581
<< polycont >>
rect -113 547 -45 581
rect 45 547 113 581
rect -34 147 34 181
rect -34 -181 34 -147
rect -113 -581 -45 -547
rect 45 -581 113 -547
<< locali >>
rect -309 685 -213 719
rect 213 685 309 719
rect -309 623 -275 685
rect 275 623 309 685
rect -129 547 -113 581
rect -45 547 -29 581
rect 29 547 45 581
rect 113 547 129 581
rect -175 488 -141 504
rect -230 285 -175 319
rect -230 223 -196 285
rect -230 -285 -196 -223
rect -17 488 17 504
rect 141 488 175 504
rect -141 285 -134 319
rect 134 285 141 319
rect 175 285 230 319
rect -50 147 -34 181
rect 34 147 50 181
rect -96 88 -62 104
rect -96 -104 -62 -88
rect 62 88 96 104
rect 62 -104 96 -88
rect -50 -181 -34 -147
rect 34 -181 50 -147
rect -230 -319 -175 -285
rect -141 -319 -134 -285
rect 134 -319 141 -285
rect -175 -504 -141 -488
rect -17 -504 17 -488
rect 196 223 230 285
rect 196 -285 230 -223
rect 175 -319 230 -285
rect 141 -504 175 -488
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 113 -581 129 -547
rect -309 -685 -275 -623
rect 275 -685 309 -623
rect -309 -719 -213 -685
rect 213 -719 309 -685
<< viali >>
rect -113 547 -45 581
rect 45 547 113 581
rect -175 331 -141 488
rect -175 273 -141 331
rect -17 331 17 488
rect -17 319 17 331
rect 141 331 175 488
rect -17 285 17 319
rect -175 -273 -141 273
rect -17 273 17 285
rect -17 197 17 273
rect -17 181 17 197
rect 141 273 175 331
rect -34 147 34 181
rect -96 -88 -62 88
rect -17 -147 17 147
rect 62 -88 96 88
rect -34 -181 34 -147
rect -175 -331 -141 -273
rect -17 -197 17 -181
rect -17 -273 17 -197
rect -17 -285 17 -273
rect 141 -273 175 273
rect -17 -319 17 -285
rect -175 -488 -141 -331
rect -17 -331 17 -319
rect -17 -488 17 -331
rect 141 -331 175 -273
rect 141 -488 175 -331
rect -113 -581 -45 -547
rect 45 -581 113 -547
<< metal1 >>
rect -125 581 -33 587
rect -125 547 -113 581
rect -45 547 -33 581
rect -125 541 -33 547
rect 33 581 125 587
rect 33 547 45 581
rect 113 547 125 581
rect 33 541 125 547
rect -181 488 -135 500
rect -181 -488 -175 488
rect -141 -488 -135 488
rect -23 488 23 500
rect -23 187 -17 488
rect -46 181 -17 187
rect 17 187 23 488
rect 135 488 181 500
rect 17 181 46 187
rect -46 147 -34 181
rect 34 147 46 181
rect -46 141 -17 147
rect -102 88 -56 100
rect -102 -88 -96 88
rect -62 -88 -56 88
rect -102 -100 -56 -88
rect -23 -141 -17 141
rect -46 -147 -17 -141
rect 17 141 46 147
rect 17 -141 23 141
rect 56 88 102 100
rect 56 -88 62 88
rect 96 -88 102 88
rect 56 -100 102 -88
rect 17 -147 46 -141
rect -46 -181 -34 -147
rect 34 -181 46 -147
rect -46 -187 -17 -181
rect -181 -500 -135 -488
rect -23 -488 -17 -187
rect 17 -187 46 -181
rect 17 -488 23 -187
rect -23 -500 23 -488
rect 135 -488 141 488
rect 175 -488 181 488
rect 135 -500 181 -488
rect -125 -547 -33 -541
rect -125 -581 -113 -547
rect -45 -581 -33 -547
rect -125 -587 -33 -581
rect 33 -547 125 -541
rect 33 -581 45 -547
rect 113 -581 125 -547
rect 33 -587 125 -581
<< properties >>
string FIXED_BBOX -213 -302 213 302
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
