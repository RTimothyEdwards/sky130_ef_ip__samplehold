magic
tech sky130A
magscale 1 2
timestamp 1718240546
<< metal3 >>
rect 2013 -17007 3394 -16918
rect 4122 -17007 7180 -16918
rect 7908 -17007 10966 -16918
rect 11694 -17007 13175 -16918
rect 2013 -18296 3394 -18207
rect 4122 -18296 7180 -18207
rect 7908 -18296 10966 -18207
rect 11694 -18296 13175 -18207
rect 2013 -19585 3394 -19496
rect 4122 -19585 7180 -19496
rect 7908 -19585 10966 -19496
rect 11694 -19585 13175 -19496
rect 2013 -20874 3394 -20785
rect 4122 -20874 7180 -20785
rect 7908 -20874 10966 -20785
rect 11694 -20874 13175 -20785
rect 2013 -22163 3394 -22074
rect 4122 -22163 7180 -22074
rect 7908 -22163 10966 -22074
rect 11694 -22163 13175 -22074
rect 2013 -23452 3395 -23363
rect 4122 -23452 7180 -23363
rect 7908 -23452 10966 -23363
rect 11694 -23452 13175 -23363
rect 2013 -24741 3394 -24652
rect 4122 -24741 7180 -24652
rect 7908 -24741 10966 -24652
rect 11694 -24741 13175 -24652
<< metal4 >>
rect 1929 -15207 13175 -15183
rect 1929 -15209 4263 -15207
rect 1929 -15526 2337 -15209
rect 3248 -15524 4263 -15209
rect 5174 -15209 8051 -15207
rect 5174 -15524 6121 -15209
rect 3248 -15526 6121 -15524
rect 7032 -15524 8051 -15209
rect 8962 -15209 11836 -15207
rect 8962 -15524 9906 -15209
rect 7032 -15526 9906 -15524
rect 10817 -15524 11836 -15209
rect 12747 -15524 13175 -15207
rect 10817 -15526 13175 -15524
rect 1929 -15549 13175 -15526
rect 1929 -15667 2025 -15549
rect 5491 -15626 5587 -15549
rect 5715 -15626 5811 -15549
rect 9277 -15667 9373 -15549
rect 9501 -15668 9597 -15549
rect 13063 -15667 13159 -15549
rect 2194 -17007 5322 -16918
rect 5980 -17007 9108 -16918
rect 9766 -17007 12894 -16918
rect 2194 -18296 5322 -18207
rect 5980 -18296 9108 -18207
rect 9766 -18296 12894 -18207
rect 2194 -19585 5322 -19496
rect 5980 -19585 9108 -19496
rect 9766 -19585 12894 -19496
rect 2194 -20874 5322 -20785
rect 5980 -20874 9108 -20785
rect 9766 -20874 12894 -20785
rect 2194 -22163 5322 -22074
rect 5980 -22163 9108 -22074
rect 9766 -22163 12894 -22074
rect 2194 -23452 5322 -23363
rect 5980 -23452 9108 -23363
rect 9766 -23452 12894 -23363
rect 2194 -24741 5322 -24652
rect 5980 -24741 9108 -24652
rect 9766 -24741 12894 -24652
<< via4 >>
rect 2337 -15526 3248 -15209
rect 4263 -15524 5174 -15207
rect 6121 -15526 7032 -15209
rect 8051 -15524 8962 -15207
rect 9906 -15526 10817 -15209
rect 11836 -15524 12747 -15207
<< metal5 >>
rect 2310 -15209 3278 -15183
rect 2310 -15526 2337 -15209
rect 3248 -15526 3278 -15209
rect 2310 -15834 3278 -15526
rect 4238 -15207 5206 -15183
rect 4238 -15524 4263 -15207
rect 5174 -15524 5206 -15207
rect 4238 -15834 5206 -15524
rect 6096 -15209 7064 -15183
rect 6096 -15526 6121 -15209
rect 7032 -15526 7064 -15209
rect 6096 -15834 7064 -15526
rect 8024 -15207 8992 -15183
rect 8024 -15524 8051 -15207
rect 8962 -15524 8992 -15207
rect 8024 -15834 8992 -15524
rect 9882 -15209 10850 -15183
rect 9882 -15526 9906 -15209
rect 10817 -15526 10850 -15209
rect 9882 -15834 10850 -15526
rect 11810 -15207 12778 -15183
rect 11810 -15524 11836 -15207
rect 12747 -15524 12778 -15207
rect 11810 -15834 12778 -15524
rect 2310 -17123 3278 -16802
rect 4238 -17123 5206 -16802
rect 6096 -17123 7064 -16802
rect 8024 -17123 8992 -16802
rect 9882 -17123 10850 -16802
rect 11810 -17123 12778 -16802
rect 2310 -18412 3278 -18091
rect 4238 -18412 5206 -18091
rect 6096 -18412 7064 -18091
rect 8024 -18412 8992 -18091
rect 9882 -18412 10850 -18091
rect 11810 -18412 12778 -18091
rect 2310 -19701 3278 -19380
rect 4238 -19701 5206 -19380
rect 6096 -19701 7064 -19380
rect 8024 -19701 8992 -19380
rect 9882 -19701 10850 -19380
rect 11810 -19701 12778 -19380
rect 2310 -20990 3278 -20669
rect 4238 -20990 5206 -20669
rect 6096 -20990 7064 -20669
rect 8024 -20990 8992 -20669
rect 9882 -20990 10850 -20669
rect 11810 -20990 12778 -20669
rect 2310 -22279 3278 -21958
rect 4238 -22279 5206 -21958
rect 6096 -22279 7064 -21958
rect 8024 -22279 8992 -21958
rect 9882 -22279 10850 -21958
rect 11810 -22279 12778 -21958
rect 2310 -23568 3278 -23247
rect 4238 -23568 5206 -23247
rect 6096 -23568 7064 -23247
rect 8024 -23568 8992 -23247
rect 9882 -23568 10850 -23247
rect 11810 -23568 12778 -23247
rect 2310 -24857 3278 -24536
rect 4238 -24857 5206 -24536
rect 6096 -24857 7064 -24536
rect 8024 -24857 8992 -24536
rect 9882 -24857 10850 -24536
rect 11810 -24857 12778 -24536
rect 3598 -26158 3918 -25920
rect 7384 -26158 7704 -25920
rect 11170 -26158 11490 -25920
rect 1997 -26553 13175 -26158
use sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt  sky130_fd_pr__cap_mim_m3_1_VCAG9S_0 paramcells
array 0 0 -1381 0 7 1289
timestamp 1718240546
transform -1 0 2744 0 1 -25341
box -650 -600 819 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt  sky130_fd_pr__cap_mim_m3_1_VCAG9S_1
array 0 0 1381 0 7 1289
timestamp 1718240546
transform 1 0 4772 0 1 -25341
box -650 -600 819 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt  sky130_fd_pr__cap_mim_m3_1_VCAG9S_2
array 0 0 -1381 0 7 1289
timestamp 1718240546
transform -1 0 6530 0 1 -25341
box -650 -600 819 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt  sky130_fd_pr__cap_mim_m3_1_VCAG9S_3
array 0 0 1381 0 7 1289
timestamp 1718240546
transform 1 0 8558 0 1 -25341
box -650 -600 819 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt  sky130_fd_pr__cap_mim_m3_1_VCAG9S_4
array 0 0 -1381 0 7 1289
timestamp 1718240546
transform -1 0 10316 0 1 -25341
box -650 -600 819 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S_alt  sky130_fd_pr__cap_mim_m3_1_VCAG9S_5
array 0 0 1381 0 7 1289
timestamp 1718240546
transform 1 0 12344 0 1 -25341
box -650 -600 819 701
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_0 paramcells
array 0 0 -1724 0 7 1289
timestamp 1718240546
transform -1 0 4471 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_1
array 0 0 1724 0 7 1289
timestamp 1718240546
transform 1 0 6831 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_2
array 0 0 -1724 0 7 1289
timestamp 1718240546
transform -1 0 8257 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_3
array 0 0 1724 0 7 1289
timestamp 1718240546
transform 1 0 10617 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_4
array 0 0 -1724 0 7 1289
timestamp 1718240546
transform -1 0 12043 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  XC2
array 0 0 1724 0 7 1289
timestamp 1718240546
transform 1 0 3045 0 1 -25341
box -851 -601 873 688
<< labels >>
flabel metal5 3731 -26364 3731 -26364 0 FreeSans 1600 0 0 0 holdval
flabel metal4 3664 -15349 3664 -15349 0 FreeSans 1600 0 0 0 vss
<< end >>
