magic
tech sky130A
magscale 1 2
timestamp 1651944383
<< metal3 >>
rect -650 10322 649 10350
rect -650 9178 565 10322
rect 629 9178 649 10322
rect -650 9150 649 9178
rect -650 9022 649 9050
rect -650 7878 565 9022
rect 629 7878 649 9022
rect -650 7850 649 7878
rect -650 7722 649 7750
rect -650 6578 565 7722
rect 629 6578 649 7722
rect -650 6550 649 6578
rect -650 6422 649 6450
rect -650 5278 565 6422
rect 629 5278 649 6422
rect -650 5250 649 5278
rect -650 5122 649 5150
rect -650 3978 565 5122
rect 629 3978 649 5122
rect -650 3950 649 3978
rect -650 3822 649 3850
rect -650 2678 565 3822
rect 629 2678 649 3822
rect -650 2650 649 2678
rect -650 2522 649 2550
rect -650 1378 565 2522
rect 629 1378 649 2522
rect -650 1350 649 1378
rect -650 1222 649 1250
rect -650 78 565 1222
rect 629 78 649 1222
rect -650 50 649 78
rect -650 -78 649 -50
rect -650 -1222 565 -78
rect 629 -1222 649 -78
rect -650 -1250 649 -1222
rect -650 -1378 649 -1350
rect -650 -2522 565 -1378
rect 629 -2522 649 -1378
rect -650 -2550 649 -2522
rect -650 -2678 649 -2650
rect -650 -3822 565 -2678
rect 629 -3822 649 -2678
rect -650 -3850 649 -3822
rect -650 -3978 649 -3950
rect -650 -5122 565 -3978
rect 629 -5122 649 -3978
rect -650 -5150 649 -5122
rect -650 -5278 649 -5250
rect -650 -6422 565 -5278
rect 629 -6422 649 -5278
rect -650 -6450 649 -6422
rect -650 -6578 649 -6550
rect -650 -7722 565 -6578
rect 629 -7722 649 -6578
rect -650 -7750 649 -7722
rect -650 -7878 649 -7850
rect -650 -9022 565 -7878
rect 629 -9022 649 -7878
rect -650 -9050 649 -9022
rect -650 -9178 649 -9150
rect -650 -10322 565 -9178
rect 629 -10322 649 -9178
rect -650 -10350 649 -10322
<< via3 >>
rect 565 9178 629 10322
rect 565 7878 629 9022
rect 565 6578 629 7722
rect 565 5278 629 6422
rect 565 3978 629 5122
rect 565 2678 629 3822
rect 565 1378 629 2522
rect 565 78 629 1222
rect 565 -1222 629 -78
rect 565 -2522 629 -1378
rect 565 -3822 629 -2678
rect 565 -5122 629 -3978
rect 565 -6422 629 -5278
rect 565 -7722 629 -6578
rect 565 -9022 629 -7878
rect 565 -10322 629 -9178
<< mimcap >>
rect -550 10210 450 10250
rect -550 9290 -510 10210
rect 410 9290 450 10210
rect -550 9250 450 9290
rect -550 8910 450 8950
rect -550 7990 -510 8910
rect 410 7990 450 8910
rect -550 7950 450 7990
rect -550 7610 450 7650
rect -550 6690 -510 7610
rect 410 6690 450 7610
rect -550 6650 450 6690
rect -550 6310 450 6350
rect -550 5390 -510 6310
rect 410 5390 450 6310
rect -550 5350 450 5390
rect -550 5010 450 5050
rect -550 4090 -510 5010
rect 410 4090 450 5010
rect -550 4050 450 4090
rect -550 3710 450 3750
rect -550 2790 -510 3710
rect 410 2790 450 3710
rect -550 2750 450 2790
rect -550 2410 450 2450
rect -550 1490 -510 2410
rect 410 1490 450 2410
rect -550 1450 450 1490
rect -550 1110 450 1150
rect -550 190 -510 1110
rect 410 190 450 1110
rect -550 150 450 190
rect -550 -190 450 -150
rect -550 -1110 -510 -190
rect 410 -1110 450 -190
rect -550 -1150 450 -1110
rect -550 -1490 450 -1450
rect -550 -2410 -510 -1490
rect 410 -2410 450 -1490
rect -550 -2450 450 -2410
rect -550 -2790 450 -2750
rect -550 -3710 -510 -2790
rect 410 -3710 450 -2790
rect -550 -3750 450 -3710
rect -550 -4090 450 -4050
rect -550 -5010 -510 -4090
rect 410 -5010 450 -4090
rect -550 -5050 450 -5010
rect -550 -5390 450 -5350
rect -550 -6310 -510 -5390
rect 410 -6310 450 -5390
rect -550 -6350 450 -6310
rect -550 -6690 450 -6650
rect -550 -7610 -510 -6690
rect 410 -7610 450 -6690
rect -550 -7650 450 -7610
rect -550 -7990 450 -7950
rect -550 -8910 -510 -7990
rect 410 -8910 450 -7990
rect -550 -8950 450 -8910
rect -550 -9290 450 -9250
rect -550 -10210 -510 -9290
rect 410 -10210 450 -9290
rect -550 -10250 450 -10210
<< mimcapcontact >>
rect -510 9290 410 10210
rect -510 7990 410 8910
rect -510 6690 410 7610
rect -510 5390 410 6310
rect -510 4090 410 5010
rect -510 2790 410 3710
rect -510 1490 410 2410
rect -510 190 410 1110
rect -510 -1110 410 -190
rect -510 -2410 410 -1490
rect -510 -3710 410 -2790
rect -510 -5010 410 -4090
rect -510 -6310 410 -5390
rect -510 -7610 410 -6690
rect -510 -8910 410 -7990
rect -510 -10210 410 -9290
<< metal4 >>
rect -102 10211 2 10400
rect 518 10338 622 10400
rect 518 10322 645 10338
rect -511 10210 411 10211
rect -511 9290 -510 10210
rect 410 9290 411 10210
rect -511 9289 411 9290
rect -102 8911 2 9289
rect 518 9178 565 10322
rect 629 9178 645 10322
rect 518 9162 645 9178
rect 518 9038 622 9162
rect 518 9022 645 9038
rect -511 8910 411 8911
rect -511 7990 -510 8910
rect 410 7990 411 8910
rect -511 7989 411 7990
rect -102 7611 2 7989
rect 518 7878 565 9022
rect 629 7878 645 9022
rect 518 7862 645 7878
rect 518 7738 622 7862
rect 518 7722 645 7738
rect -511 7610 411 7611
rect -511 6690 -510 7610
rect 410 6690 411 7610
rect -511 6689 411 6690
rect -102 6311 2 6689
rect 518 6578 565 7722
rect 629 6578 645 7722
rect 518 6562 645 6578
rect 518 6438 622 6562
rect 518 6422 645 6438
rect -511 6310 411 6311
rect -511 5390 -510 6310
rect 410 5390 411 6310
rect -511 5389 411 5390
rect -102 5011 2 5389
rect 518 5278 565 6422
rect 629 5278 645 6422
rect 518 5262 645 5278
rect 518 5138 622 5262
rect 518 5122 645 5138
rect -511 5010 411 5011
rect -511 4090 -510 5010
rect 410 4090 411 5010
rect -511 4089 411 4090
rect -102 3711 2 4089
rect 518 3978 565 5122
rect 629 3978 645 5122
rect 518 3962 645 3978
rect 518 3838 622 3962
rect 518 3822 645 3838
rect -511 3710 411 3711
rect -511 2790 -510 3710
rect 410 2790 411 3710
rect -511 2789 411 2790
rect -102 2411 2 2789
rect 518 2678 565 3822
rect 629 2678 645 3822
rect 518 2662 645 2678
rect 518 2538 622 2662
rect 518 2522 645 2538
rect -511 2410 411 2411
rect -511 1490 -510 2410
rect 410 1490 411 2410
rect -511 1489 411 1490
rect -102 1111 2 1489
rect 518 1378 565 2522
rect 629 1378 645 2522
rect 518 1362 645 1378
rect 518 1238 622 1362
rect 518 1222 645 1238
rect -511 1110 411 1111
rect -511 190 -510 1110
rect 410 190 411 1110
rect -511 189 411 190
rect -102 -189 2 189
rect 518 78 565 1222
rect 629 78 645 1222
rect 518 62 645 78
rect 518 -62 622 62
rect 518 -78 645 -62
rect -511 -190 411 -189
rect -511 -1110 -510 -190
rect 410 -1110 411 -190
rect -511 -1111 411 -1110
rect -102 -1489 2 -1111
rect 518 -1222 565 -78
rect 629 -1222 645 -78
rect 518 -1238 645 -1222
rect 518 -1362 622 -1238
rect 518 -1378 645 -1362
rect -511 -1490 411 -1489
rect -511 -2410 -510 -1490
rect 410 -2410 411 -1490
rect -511 -2411 411 -2410
rect -102 -2789 2 -2411
rect 518 -2522 565 -1378
rect 629 -2522 645 -1378
rect 518 -2538 645 -2522
rect 518 -2662 622 -2538
rect 518 -2678 645 -2662
rect -511 -2790 411 -2789
rect -511 -3710 -510 -2790
rect 410 -3710 411 -2790
rect -511 -3711 411 -3710
rect -102 -4089 2 -3711
rect 518 -3822 565 -2678
rect 629 -3822 645 -2678
rect 518 -3838 645 -3822
rect 518 -3962 622 -3838
rect 518 -3978 645 -3962
rect -511 -4090 411 -4089
rect -511 -5010 -510 -4090
rect 410 -5010 411 -4090
rect -511 -5011 411 -5010
rect -102 -5389 2 -5011
rect 518 -5122 565 -3978
rect 629 -5122 645 -3978
rect 518 -5138 645 -5122
rect 518 -5262 622 -5138
rect 518 -5278 645 -5262
rect -511 -5390 411 -5389
rect -511 -6310 -510 -5390
rect 410 -6310 411 -5390
rect -511 -6311 411 -6310
rect -102 -6689 2 -6311
rect 518 -6422 565 -5278
rect 629 -6422 645 -5278
rect 518 -6438 645 -6422
rect 518 -6562 622 -6438
rect 518 -6578 645 -6562
rect -511 -6690 411 -6689
rect -511 -7610 -510 -6690
rect 410 -7610 411 -6690
rect -511 -7611 411 -7610
rect -102 -7989 2 -7611
rect 518 -7722 565 -6578
rect 629 -7722 645 -6578
rect 518 -7738 645 -7722
rect 518 -7862 622 -7738
rect 518 -7878 645 -7862
rect -511 -7990 411 -7989
rect -511 -8910 -510 -7990
rect 410 -8910 411 -7990
rect -511 -8911 411 -8910
rect -102 -9289 2 -8911
rect 518 -9022 565 -7878
rect 629 -9022 645 -7878
rect 518 -9038 645 -9022
rect 518 -9162 622 -9038
rect 518 -9178 645 -9162
rect -511 -9290 411 -9289
rect -511 -10210 -510 -9290
rect 410 -10210 411 -9290
rect -511 -10211 411 -10210
rect -102 -10400 2 -10211
rect 518 -10322 565 -9178
rect 629 -10322 645 -9178
rect 518 -10338 645 -10322
rect 518 -10400 622 -10338
<< properties >>
string FIXED_BBOX -650 9150 550 10350
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.0 l 5.0 val 53.8 carea 2.00 cperi 0.19 nx 1 ny 16 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
