magic
tech sky130A
magscale 1 2
timestamp 1717691772
<< pwell >>
rect -782 -1832 782 1832
<< psubdiff >>
rect -746 1762 -650 1796
rect 650 1762 746 1796
rect -746 1700 -712 1762
rect 712 1700 746 1762
rect -746 -1762 -712 -1700
rect 712 -1762 746 -1700
rect -746 -1796 -650 -1762
rect 650 -1796 746 -1762
<< psubdiffcont >>
rect -650 1762 650 1796
rect -746 -1700 -712 1700
rect 712 -1700 746 1700
rect -650 -1796 650 -1762
<< xpolycontact >>
rect -616 1234 -546 1666
rect -616 -1666 -546 -1234
rect -450 1234 -380 1666
rect -450 -1666 -380 -1234
rect -284 1234 -214 1666
rect -284 -1666 -214 -1234
rect -118 1234 -48 1666
rect -118 -1666 -48 -1234
rect 48 1234 118 1666
rect 48 -1666 118 -1234
rect 214 1234 284 1666
rect 214 -1666 284 -1234
rect 380 1234 450 1666
rect 380 -1666 450 -1234
rect 546 1234 616 1666
rect 546 -1666 616 -1234
<< xpolyres >>
rect -616 -1234 -546 1234
rect -450 -1234 -380 1234
rect -284 -1234 -214 1234
rect -118 -1234 -48 1234
rect 48 -1234 118 1234
rect 214 -1234 284 1234
rect 380 -1234 450 1234
rect 546 -1234 616 1234
<< locali >>
rect -746 1762 -650 1796
rect 650 1762 746 1796
rect -746 1700 -712 1762
rect 712 1700 746 1762
rect -746 -1762 -712 -1700
rect 712 -1762 746 -1700
rect -746 -1796 -650 -1762
rect 650 -1796 746 -1762
<< viali >>
rect -600 1251 -562 1648
rect -434 1251 -396 1648
rect -268 1251 -230 1648
rect -102 1251 -64 1648
rect 64 1251 102 1648
rect 230 1251 268 1648
rect 396 1251 434 1648
rect 562 1251 600 1648
rect -600 -1648 -562 -1251
rect -434 -1648 -396 -1251
rect -268 -1648 -230 -1251
rect -102 -1648 -64 -1251
rect 64 -1648 102 -1251
rect 230 -1648 268 -1251
rect 396 -1648 434 -1251
rect 562 -1648 600 -1251
<< metal1 >>
rect -606 1648 -556 1660
rect -606 1251 -600 1648
rect -562 1251 -556 1648
rect -606 1239 -556 1251
rect -440 1648 -390 1660
rect -440 1251 -434 1648
rect -396 1251 -390 1648
rect -440 1239 -390 1251
rect -274 1648 -224 1660
rect -274 1251 -268 1648
rect -230 1251 -224 1648
rect -274 1239 -224 1251
rect -108 1648 -58 1660
rect -108 1251 -102 1648
rect -64 1251 -58 1648
rect -108 1239 -58 1251
rect 58 1648 108 1660
rect 58 1251 64 1648
rect 102 1251 108 1648
rect 58 1239 108 1251
rect 224 1648 274 1660
rect 224 1251 230 1648
rect 268 1251 274 1648
rect 224 1239 274 1251
rect 390 1648 440 1660
rect 390 1251 396 1648
rect 434 1251 440 1648
rect 390 1239 440 1251
rect 556 1648 606 1660
rect 556 1251 562 1648
rect 600 1251 606 1648
rect 556 1239 606 1251
rect -606 -1251 -556 -1239
rect -606 -1648 -600 -1251
rect -562 -1648 -556 -1251
rect -606 -1660 -556 -1648
rect -440 -1251 -390 -1239
rect -440 -1648 -434 -1251
rect -396 -1648 -390 -1251
rect -440 -1660 -390 -1648
rect -274 -1251 -224 -1239
rect -274 -1648 -268 -1251
rect -230 -1648 -224 -1251
rect -274 -1660 -224 -1648
rect -108 -1251 -58 -1239
rect -108 -1648 -102 -1251
rect -64 -1648 -58 -1251
rect -108 -1660 -58 -1648
rect 58 -1251 108 -1239
rect 58 -1648 64 -1251
rect 102 -1648 108 -1251
rect 58 -1660 108 -1648
rect 224 -1251 274 -1239
rect 224 -1648 230 -1251
rect 268 -1648 274 -1251
rect 224 -1660 274 -1648
rect 390 -1251 440 -1239
rect 390 -1648 396 -1251
rect 434 -1648 440 -1251
rect 390 -1660 440 -1648
rect 556 -1251 606 -1239
rect 556 -1648 562 -1251
rect 600 -1648 606 -1251
rect 556 -1660 606 -1648
<< properties >>
string FIXED_BBOX -729 -1779 729 1779
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 12.5 m 1 nx 8 wmin 0.350 lmin 0.50 rho 2000 val 72.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
