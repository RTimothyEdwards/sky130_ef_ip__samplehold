magic
tech sky130A
magscale 1 2
timestamp 1717692607
<< pwell >>
rect -437 -358 437 358
<< mvnnmos >>
rect -209 -100 -29 100
rect 29 -100 209 100
<< mvndiff >>
rect -267 88 -209 100
rect -267 -88 -255 88
rect -221 -88 -209 88
rect -267 -100 -209 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 209 88 267 100
rect 209 -88 221 88
rect 255 -88 267 88
rect 209 -100 267 -88
<< mvndiffc >>
rect -255 -88 -221 88
rect -17 -88 17 88
rect 221 -88 255 88
<< mvpsubdiff >>
rect -401 310 401 322
rect -401 276 -293 310
rect 293 276 401 310
rect -401 264 401 276
rect -401 214 -343 264
rect -401 -214 -389 214
rect -355 -214 -343 214
rect -401 -264 -343 -214
rect 343 -264 401 264
rect -401 -276 401 -264
rect -401 -310 -293 -276
rect 293 -310 401 -276
rect -401 -322 401 -310
<< mvpsubdiffcont >>
rect -293 276 293 310
rect -389 -214 -355 214
rect -293 -310 293 -276
<< poly >>
rect -209 172 -29 188
rect -209 138 -193 172
rect -45 138 -29 172
rect -209 100 -29 138
rect 29 172 209 188
rect 29 138 45 172
rect 193 138 209 172
rect 29 100 209 138
rect -209 -138 -29 -100
rect -209 -172 -193 -138
rect -45 -172 -29 -138
rect -209 -188 -29 -172
rect 29 -138 209 -100
rect 29 -172 45 -138
rect 193 -172 209 -138
rect 29 -188 209 -172
<< polycont >>
rect -193 138 -45 172
rect 45 138 193 172
rect -193 -172 -45 -138
rect 45 -172 193 -138
<< locali >>
rect -389 276 -293 310
rect 293 276 389 310
rect -389 214 -355 276
rect -209 138 -193 172
rect -45 138 -29 172
rect 29 138 45 172
rect 193 138 209 172
rect -255 88 -221 104
rect -255 -104 -221 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 221 88 255 104
rect 221 -104 255 -88
rect -209 -172 -193 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 193 -172 209 -138
rect -389 -276 -355 -214
rect 355 -276 389 276
rect -389 -310 -293 -276
rect 293 -310 389 -276
<< viali >>
rect -193 138 -45 172
rect 45 138 193 172
rect -255 -88 -221 88
rect -17 -88 17 88
rect 221 -88 255 88
rect -193 -172 -45 -138
rect 45 -172 193 -138
<< metal1 >>
rect -205 172 -33 178
rect -205 138 -193 172
rect -45 138 -33 172
rect -205 132 -33 138
rect 33 172 205 178
rect 33 138 45 172
rect 193 138 205 172
rect 33 132 205 138
rect -261 88 -215 100
rect -261 -88 -255 88
rect -221 -88 -215 88
rect -261 -100 -215 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 215 88 261 100
rect 215 -88 221 88
rect 255 -88 261 88
rect 215 -100 261 -88
rect -205 -138 -33 -132
rect -205 -172 -193 -138
rect -45 -172 -33 -138
rect -205 -178 -33 -172
rect 33 -138 205 -132
rect 33 -172 45 -138
rect 193 -172 205 -138
rect 33 -178 205 -172
<< properties >>
string FIXED_BBOX -372 -293 372 293
string gencell sky130_fd_pr__nfet_05v0_nvt
string library sky130
string parameters w 1.0 l 0.9 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.90 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
