magic
tech sky130A
timestamp 1718240546
<< metal1 >>
rect 7974 -3963 7977 -3937
rect 8108 -3963 8111 -3937
<< via1 >>
rect 7977 -3963 8108 -3937
<< metal2 >>
rect 7977 -3937 8108 -3934
rect 7977 -3966 8108 -3963
<< end >>
