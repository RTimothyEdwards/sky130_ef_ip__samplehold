magic
tech sky130A
magscale 1 2
timestamp 1718240546
<< nwell >>
rect -466 -397 466 397
<< mvpmos >>
rect -208 -100 -108 100
rect -50 -100 50 100
rect 108 -100 208 100
<< mvpdiff >>
rect -266 88 -208 100
rect -266 -88 -254 88
rect -220 -88 -208 88
rect -266 -100 -208 -88
rect -108 88 -50 100
rect -108 -88 -96 88
rect -62 -88 -50 88
rect -108 -100 -50 -88
rect 50 88 108 100
rect 50 -88 62 88
rect 96 -88 108 88
rect 50 -100 108 -88
rect 208 88 266 100
rect 208 -88 220 88
rect 254 -88 266 88
rect 208 -100 266 -88
<< mvpdiffc >>
rect -254 -88 -220 88
rect -96 -88 -62 88
rect 62 -88 96 88
rect 220 -88 254 88
<< mvnsubdiff >>
rect -400 319 400 331
rect -400 285 -292 319
rect 292 285 400 319
rect -400 273 400 285
rect -400 223 -342 273
rect -400 -223 -388 223
rect -354 -223 -342 223
rect 342 223 400 273
rect -400 -273 -342 -223
rect 342 -223 354 223
rect 388 -223 400 223
rect 342 -273 400 -223
rect -400 -285 400 -273
rect -400 -319 -292 -285
rect 292 -319 400 -285
rect -400 -331 400 -319
<< mvnsubdiffcont >>
rect -292 285 292 319
rect -388 -223 -354 223
rect 354 -223 388 223
rect -292 -319 292 -285
<< poly >>
rect -208 181 -108 197
rect -208 147 -192 181
rect -124 147 -108 181
rect -208 100 -108 147
rect -50 181 50 197
rect -50 147 -34 181
rect 34 147 50 181
rect -50 100 50 147
rect 108 181 208 197
rect 108 147 124 181
rect 192 147 208 181
rect 108 100 208 147
rect -208 -147 -108 -100
rect -208 -181 -192 -147
rect -124 -181 -108 -147
rect -208 -197 -108 -181
rect -50 -147 50 -100
rect -50 -181 -34 -147
rect 34 -181 50 -147
rect -50 -197 50 -181
rect 108 -147 208 -100
rect 108 -181 124 -147
rect 192 -181 208 -147
rect 108 -197 208 -181
<< polycont >>
rect -192 147 -124 181
rect -34 147 34 181
rect 124 147 192 181
rect -192 -181 -124 -147
rect -34 -181 34 -147
rect 124 -181 192 -147
<< locali >>
rect -388 285 -292 319
rect 292 285 388 319
rect -388 223 -354 285
rect 354 223 388 285
rect -208 147 -192 181
rect -124 147 -108 181
rect -50 147 -34 181
rect 34 147 50 181
rect 108 147 124 181
rect 192 147 208 181
rect -254 88 -220 104
rect -254 -104 -220 -88
rect -96 88 -62 104
rect -96 -104 -62 -88
rect 62 88 96 104
rect 62 -104 96 -88
rect 220 88 254 104
rect 220 -104 254 -88
rect -208 -181 -192 -147
rect -124 -181 -108 -147
rect -50 -181 -34 -147
rect 34 -181 50 -147
rect 108 -181 124 -147
rect 192 -181 208 -147
rect -388 -285 -354 -223
rect 354 -285 388 -223
rect -388 -319 -292 -285
rect 292 -319 388 -285
<< viali >>
rect -192 147 -124 181
rect -34 147 34 181
rect 124 147 192 181
rect -254 -88 -220 88
rect -96 -88 -62 88
rect 62 -88 96 88
rect 220 -88 254 88
rect -192 -181 -124 -147
rect -34 -181 34 -147
rect 124 -181 192 -147
<< metal1 >>
rect -204 181 -112 187
rect -204 147 -192 181
rect -124 147 -112 181
rect -204 141 -112 147
rect -46 181 46 187
rect -46 147 -34 181
rect 34 147 46 181
rect -46 141 46 147
rect 112 181 204 187
rect 112 147 124 181
rect 192 147 204 181
rect 112 141 204 147
rect -260 88 -214 100
rect -260 -88 -254 88
rect -220 -88 -214 88
rect -260 -100 -214 -88
rect -102 88 -56 100
rect -102 -88 -96 88
rect -62 -88 -56 88
rect -102 -100 -56 -88
rect 56 88 102 100
rect 56 -88 62 88
rect 96 -88 102 88
rect 56 -100 102 -88
rect 214 88 260 100
rect 214 -88 220 88
rect 254 -88 260 88
rect 214 -100 260 -88
rect -204 -147 -112 -141
rect -204 -181 -192 -147
rect -124 -181 -112 -147
rect -204 -187 -112 -181
rect -46 -147 46 -141
rect -46 -181 -34 -147
rect 34 -181 46 -147
rect -46 -187 46 -181
rect 112 -147 204 -141
rect 112 -181 124 -147
rect 192 -181 204 -147
rect 112 -187 204 -181
<< properties >>
string FIXED_BBOX -371 -302 371 302
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
