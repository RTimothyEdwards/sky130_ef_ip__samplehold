magic
tech sky130A
magscale 1 2
timestamp 1717690002
<< nwell >>
rect -308 -397 308 397
<< mvpmos >>
rect -50 -100 50 100
<< mvpdiff >>
rect -108 88 -50 100
rect -108 -88 -96 88
rect -62 -88 -50 88
rect -108 -100 -50 -88
rect 50 88 108 100
rect 50 -88 62 88
rect 96 -88 108 88
rect 50 -100 108 -88
<< mvpdiffc >>
rect -96 -88 -62 88
rect 62 -88 96 88
<< mvnsubdiff >>
rect -242 319 242 331
rect -242 285 -134 319
rect 134 285 242 319
rect -242 273 242 285
rect -242 223 -184 273
rect -242 -223 -230 223
rect -196 -223 -184 223
rect 184 223 242 273
rect -242 -273 -184 -223
rect 184 -223 196 223
rect 230 -223 242 223
rect 184 -273 242 -223
rect -242 -285 242 -273
rect -242 -319 -134 -285
rect 134 -319 242 -285
rect -242 -331 242 -319
<< mvnsubdiffcont >>
rect -134 285 134 319
rect -230 -223 -196 223
rect 196 -223 230 223
rect -134 -319 134 -285
<< poly >>
rect -50 181 50 197
rect -50 147 -34 181
rect 34 147 50 181
rect -50 100 50 147
rect -50 -147 50 -100
rect -50 -181 -34 -147
rect 34 -181 50 -147
rect -50 -197 50 -181
<< polycont >>
rect -34 147 34 181
rect -34 -181 34 -147
<< locali >>
rect -230 285 -134 319
rect 134 285 230 319
rect -230 223 -196 285
rect 196 223 230 285
rect -50 147 -34 181
rect 34 147 50 181
rect -96 88 -62 104
rect -96 -104 -62 -88
rect 62 88 96 104
rect 62 -104 96 -88
rect -50 -181 -34 -147
rect 34 -181 50 -147
rect -230 -285 -196 -223
rect 196 -285 230 -223
rect -230 -319 -134 -285
rect 134 -319 230 -285
<< viali >>
rect -34 147 34 181
rect -96 -88 -62 88
rect 62 -88 96 88
rect -34 -181 34 -147
<< metal1 >>
rect -46 181 46 187
rect -46 147 -34 181
rect 34 147 46 181
rect -46 141 46 147
rect -102 88 -56 100
rect -102 -88 -96 88
rect -62 -88 -56 88
rect -102 -100 -56 -88
rect 56 88 102 100
rect 56 -88 62 88
rect 96 -88 102 88
rect 56 -100 102 -88
rect -46 -147 46 -141
rect -46 -181 -34 -147
rect 34 -181 46 -147
rect -46 -187 46 -181
<< properties >>
string FIXED_BBOX -213 -302 213 302
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
