magic
tech sky130A
magscale 1 2
timestamp 1718228583
<< dnwell >>
rect 229 230 4145 10887
<< nwell >>
rect 120 10681 4254 10996
rect 120 436 435 10681
rect 3939 436 4254 10681
rect 120 121 4254 436
<< mvpsubdiff >>
rect 0 11093 60 11127
rect 4316 11093 4376 11127
rect 0 11067 34 11093
rect 4342 11067 4376 11093
rect 0 34 34 130
rect 4342 34 4376 130
rect 0 0 60 34
rect 4316 0 4376 34
<< mvnsubdiff >>
rect 186 10910 4188 10930
rect 186 10876 266 10910
rect 4108 10876 4188 10910
rect 186 10856 4188 10876
rect 186 10850 260 10856
rect 186 267 206 10850
rect 240 267 260 10850
rect 186 261 260 267
rect 4114 10850 4188 10856
rect 4114 267 4134 10850
rect 4168 267 4188 10850
rect 4114 261 4188 267
rect 186 241 4188 261
rect 186 207 266 241
rect 4108 207 4188 241
rect 186 187 4188 207
<< mvpsubdiffcont >>
rect 60 11093 4316 11127
rect 0 130 34 11067
rect 4342 130 4376 11067
rect 60 0 4316 34
<< mvnsubdiffcont >>
rect 266 10876 4108 10910
rect 206 267 240 10850
rect 4134 267 4168 10850
rect 266 207 4108 241
<< locali >>
rect 0 11127 4377 11129
rect 0 11093 60 11127
rect 4316 11093 4377 11127
rect 0 11071 164 11093
rect 0 11067 45 11071
rect 34 211 45 11067
rect 89 11049 164 11071
rect 4228 11078 4377 11093
rect 4228 11049 4301 11078
rect 4347 11067 4377 11078
rect 89 11029 4301 11049
rect 89 211 108 11029
rect 34 130 108 211
rect 179 10939 283 10943
rect 179 10920 4188 10939
rect 179 10910 281 10920
rect 4083 10910 4188 10920
rect 179 10876 266 10910
rect 4108 10876 4188 10910
rect 179 10868 281 10876
rect 4083 10868 4188 10876
rect 179 10850 4188 10868
rect 179 10840 206 10850
rect 240 10848 4134 10850
rect 240 10840 283 10848
rect 179 292 202 10840
rect 247 292 283 10840
rect 4087 10827 4134 10848
rect 372 10706 3973 10732
rect 372 10671 521 10706
rect 3770 10703 3973 10706
rect 3770 10671 3930 10703
rect 372 10643 3930 10671
rect 372 10410 542 10643
rect 372 3817 383 10410
rect 437 4472 542 10410
rect 3884 4472 3930 10643
rect 437 4440 3930 4472
rect 437 4398 646 4440
rect 3790 4398 3930 4440
rect 437 4371 3930 4398
rect 437 3857 542 4371
rect 3884 3857 3930 4371
rect 437 3841 3930 3857
rect 437 3817 677 3841
rect 372 3806 677 3817
rect 2924 3839 3930 3841
rect 2924 3806 3114 3839
rect 372 3805 3114 3806
rect 3806 3805 3930 3839
rect 372 3768 3930 3805
rect 427 3666 3930 3696
rect 427 3665 2232 3666
rect 427 3617 475 3665
rect 2008 3619 2232 3665
rect 2946 3662 3930 3666
rect 2946 3619 3123 3662
rect 2008 3617 3123 3619
rect 427 3615 3123 3617
rect 3799 3615 3930 3662
rect 427 3585 3930 3615
rect 448 3090 559 3585
rect 3880 3128 3930 3585
rect 3969 3768 3973 10703
rect 3969 3695 3979 3696
rect 3969 3128 3991 3695
rect 3880 3090 3991 3128
rect 439 2979 3991 3090
rect 4087 3082 4124 10827
rect 4087 3055 4134 3082
rect 595 2804 3905 2827
rect 595 2719 3824 2804
rect 595 2251 703 2719
rect 3797 2251 3824 2719
rect 594 2221 3824 2251
rect 594 2170 864 2221
rect 2214 2196 3824 2221
rect 3879 2196 3905 2804
rect 2214 2170 3905 2196
rect 594 2143 3905 2170
rect 1193 2028 3905 2032
rect 586 2000 3905 2028
rect 586 1963 734 2000
rect 2742 1987 3905 2000
rect 2742 1963 3825 1987
rect 586 1947 3825 1963
rect 586 1448 687 1947
rect 893 1923 3825 1947
rect 893 1508 935 1923
rect 892 1448 935 1508
rect 586 1443 935 1448
rect 973 1918 3825 1923
rect 973 1910 1193 1918
rect 973 1443 1110 1910
rect 586 1442 1110 1443
rect 1151 1448 1193 1910
rect 2526 1448 2654 1786
rect 3791 1448 3825 1918
rect 1151 1442 3825 1448
rect 586 1419 3825 1442
rect 586 1371 1297 1419
rect 2190 1379 3825 1419
rect 3880 1379 3905 1987
rect 2190 1371 3905 1379
rect 586 1334 3905 1371
rect 892 1203 1193 1334
rect 442 1183 4015 1203
rect 442 1169 3960 1183
rect 442 1133 564 1169
rect 3290 1133 3960 1169
rect 442 1095 3960 1133
rect 442 742 537 1095
rect 442 597 459 742
rect 506 597 537 742
rect 442 548 537 597
rect 3881 548 3960 1095
rect 442 519 3960 548
rect 4000 519 4015 1183
rect 442 516 4015 519
rect 442 479 454 516
rect 3919 479 4015 516
rect 442 442 4015 479
rect 179 267 206 292
rect 240 281 283 292
rect 240 267 4134 281
rect 4168 3055 4188 10850
rect 4168 267 4195 281
rect 179 253 4195 267
rect 179 199 255 253
rect 4117 199 4195 253
rect 179 169 4195 199
rect 0 102 108 130
rect 4278 102 4301 11029
rect 4376 130 4377 11067
rect 0 72 4301 102
rect 0 34 148 72
rect 4259 70 4301 72
rect 4347 70 4377 130
rect 4259 34 4377 70
rect 0 0 60 34
rect 4316 0 4377 34
<< viali >>
rect 164 11093 4228 11095
rect 45 211 89 11071
rect 164 11049 4228 11093
rect 4301 11067 4347 11078
rect 281 10910 4083 10920
rect 281 10876 4083 10910
rect 281 10868 4083 10876
rect 202 292 206 10840
rect 206 292 240 10840
rect 240 292 247 10840
rect 521 10671 3770 10706
rect 383 3817 437 10410
rect 646 4398 3790 4440
rect 677 3806 2924 3841
rect 3114 3805 3806 3839
rect 475 3617 2008 3665
rect 2232 3619 2946 3666
rect 3123 3615 3799 3662
rect 3930 3128 3969 10703
rect 4124 3082 4134 10827
rect 4134 3082 4167 10827
rect 864 2170 2214 2221
rect 3824 2196 3879 2804
rect 734 1963 2742 2000
rect 935 1443 973 1923
rect 1110 1442 1151 1910
rect 1297 1371 2190 1419
rect 3825 1379 3880 1987
rect 564 1133 3290 1169
rect 459 597 506 742
rect 3960 519 4000 1183
rect 454 479 3919 516
rect 255 241 4117 253
rect 255 207 266 241
rect 266 207 4108 241
rect 4108 207 4117 241
rect 255 199 4117 207
rect 4301 130 4342 11067
rect 4342 130 4347 11067
rect 148 34 4259 72
rect 4301 70 4347 130
rect 148 26 4259 34
<< metal1 >>
rect 0 11095 4377 11129
rect 0 11071 164 11095
rect 0 211 45 11071
rect 89 11049 164 11071
rect 4228 11078 4377 11095
rect 4228 11049 4301 11078
rect 89 11029 4301 11049
rect 89 211 108 11029
rect 0 102 108 211
rect 179 10939 283 10943
rect 179 10920 4188 10939
rect 179 10868 281 10920
rect 4083 10868 4188 10920
rect 179 10848 4188 10868
rect 179 10840 283 10848
rect 179 292 202 10840
rect 247 4493 283 10840
rect 353 10733 458 10848
rect 3907 10734 4012 10848
rect 4087 10827 4188 10848
rect 3907 10733 4014 10734
rect 353 10732 4014 10733
rect 350 10718 4014 10732
rect 350 10706 544 10718
rect 3758 10706 4014 10718
rect 350 10671 521 10706
rect 3770 10703 4014 10706
rect 3770 10671 3930 10703
rect 350 10664 544 10671
rect 3758 10664 3930 10671
rect 350 10644 3930 10664
rect 350 10428 457 10644
rect 350 4493 360 10428
rect 247 4375 360 4493
rect 247 3693 283 4375
rect 350 3693 360 4375
rect 247 3584 360 3693
rect 247 292 283 3584
rect 350 3385 360 3584
rect 446 3671 457 10428
rect 505 10568 671 10572
rect 850 10568 882 10572
rect 1008 10568 1040 10572
rect 1166 10568 1198 10572
rect 1324 10568 1356 10572
rect 1482 10568 1514 10572
rect 1640 10568 1672 10572
rect 1798 10568 1830 10572
rect 1956 10568 1988 10572
rect 2114 10568 2146 10572
rect 2272 10568 2304 10572
rect 2430 10568 2462 10572
rect 2588 10568 2620 10572
rect 2746 10568 2778 10572
rect 2904 10568 2936 10572
rect 3062 10568 3094 10572
rect 3220 10568 3252 10572
rect 3378 10568 3410 10572
rect 3536 10568 3568 10572
rect 3694 10568 3726 10572
rect 505 10531 3765 10568
rect 505 10526 671 10531
rect 505 10244 552 10526
rect 505 10240 671 10244
rect 692 10240 724 10531
rect 850 10240 882 10531
rect 1008 10240 1040 10531
rect 1166 10240 1198 10531
rect 1324 10240 1356 10531
rect 1482 10240 1514 10531
rect 1640 10240 1672 10531
rect 1798 10240 1830 10531
rect 1956 10240 1988 10531
rect 2114 10240 2146 10531
rect 2272 10240 2304 10531
rect 2430 10240 2462 10531
rect 2588 10240 2620 10531
rect 2746 10240 2778 10531
rect 2904 10240 2936 10531
rect 3062 10240 3094 10531
rect 3220 10240 3252 10531
rect 3378 10240 3410 10531
rect 3536 10240 3568 10531
rect 3694 10240 3726 10531
rect 505 10203 3757 10240
rect 505 10198 671 10203
rect 505 10136 552 10198
rect 505 10132 671 10136
rect 692 10132 724 10203
rect 850 10132 882 10203
rect 1008 10132 1040 10203
rect 1166 10132 1198 10203
rect 1324 10132 1356 10203
rect 1482 10132 1514 10203
rect 1640 10132 1672 10203
rect 1798 10132 1830 10203
rect 1956 10132 1988 10203
rect 2114 10132 2146 10203
rect 2272 10132 2304 10203
rect 2430 10132 2462 10203
rect 2588 10132 2620 10203
rect 2746 10132 2778 10203
rect 2904 10132 2936 10203
rect 3062 10132 3094 10203
rect 3220 10132 3252 10203
rect 3378 10132 3410 10203
rect 3536 10132 3568 10203
rect 3694 10132 3726 10203
rect 505 10095 3765 10132
rect 505 10090 671 10095
rect 505 9808 552 10090
rect 505 9804 671 9808
rect 692 9804 724 10095
rect 850 9804 882 10095
rect 1008 9804 1040 10095
rect 1166 9804 1198 10095
rect 1324 9804 1356 10095
rect 1482 9804 1514 10095
rect 1640 9804 1672 10095
rect 1798 9804 1830 10095
rect 1956 9804 1988 10095
rect 2114 9804 2146 10095
rect 2272 9804 2304 10095
rect 2430 9804 2462 10095
rect 2588 9804 2620 10095
rect 2746 9804 2778 10095
rect 2904 9804 2936 10095
rect 3062 9804 3094 10095
rect 3220 9804 3252 10095
rect 3378 9804 3410 10095
rect 3536 9804 3568 10095
rect 3694 9804 3726 10095
rect 505 9767 3757 9804
rect 505 9762 671 9767
rect 505 9700 552 9762
rect 505 9696 671 9700
rect 692 9696 724 9767
rect 850 9696 882 9767
rect 1008 9696 1040 9767
rect 1166 9696 1198 9767
rect 1324 9696 1356 9767
rect 1482 9696 1514 9767
rect 1640 9696 1672 9767
rect 1798 9696 1830 9767
rect 1956 9696 1988 9767
rect 2114 9696 2146 9767
rect 2272 9696 2304 9767
rect 2430 9696 2462 9767
rect 2588 9696 2620 9767
rect 2746 9696 2778 9767
rect 2904 9696 2936 9767
rect 3062 9696 3094 9767
rect 3220 9696 3252 9767
rect 3378 9696 3410 9767
rect 3536 9696 3568 9767
rect 3694 9696 3726 9767
rect 505 9659 3765 9696
rect 505 9654 671 9659
rect 505 9372 552 9654
rect 505 9368 671 9372
rect 692 9368 724 9659
rect 850 9368 882 9659
rect 1008 9368 1040 9659
rect 1166 9368 1198 9659
rect 1324 9368 1356 9659
rect 1482 9368 1514 9659
rect 1640 9368 1672 9659
rect 1798 9368 1830 9659
rect 1956 9368 1988 9659
rect 2114 9368 2146 9659
rect 2272 9368 2304 9659
rect 2430 9368 2462 9659
rect 2588 9368 2620 9659
rect 2746 9368 2778 9659
rect 2904 9368 2936 9659
rect 3062 9368 3094 9659
rect 3220 9368 3252 9659
rect 3378 9368 3410 9659
rect 3536 9368 3568 9659
rect 3694 9368 3726 9659
rect 505 9331 3757 9368
rect 505 9326 671 9331
rect 505 9264 552 9326
rect 505 9260 671 9264
rect 692 9260 724 9331
rect 850 9260 882 9331
rect 1008 9260 1040 9331
rect 1166 9260 1198 9331
rect 1324 9260 1356 9331
rect 1482 9260 1514 9331
rect 1640 9260 1672 9331
rect 1798 9260 1830 9331
rect 1956 9260 1988 9331
rect 2114 9260 2146 9331
rect 2272 9260 2304 9331
rect 2430 9260 2462 9331
rect 2588 9260 2620 9331
rect 2746 9260 2778 9331
rect 2904 9260 2936 9331
rect 3062 9260 3094 9331
rect 3220 9260 3252 9331
rect 3378 9260 3410 9331
rect 3536 9260 3568 9331
rect 3694 9260 3726 9331
rect 505 9223 3765 9260
rect 505 9218 671 9223
rect 505 8936 552 9218
rect 505 8932 671 8936
rect 692 8932 724 9223
rect 850 8932 882 9223
rect 1008 8932 1040 9223
rect 1166 8932 1198 9223
rect 1324 8932 1356 9223
rect 1482 8932 1514 9223
rect 1640 8932 1672 9223
rect 1798 8932 1830 9223
rect 1956 8932 1988 9223
rect 2114 8932 2146 9223
rect 2272 8932 2304 9223
rect 2430 8932 2462 9223
rect 2588 8932 2620 9223
rect 2746 8932 2778 9223
rect 2904 8932 2936 9223
rect 3062 8932 3094 9223
rect 3220 8932 3252 9223
rect 3378 8932 3410 9223
rect 3536 8932 3568 9223
rect 3694 8932 3726 9223
rect 505 8895 3757 8932
rect 505 8890 671 8895
rect 505 8828 552 8890
rect 505 8824 671 8828
rect 692 8824 724 8895
rect 850 8824 882 8895
rect 1008 8824 1040 8895
rect 1166 8824 1198 8895
rect 1324 8824 1356 8895
rect 1482 8824 1514 8895
rect 1640 8824 1672 8895
rect 1798 8824 1830 8895
rect 1956 8824 1988 8895
rect 2114 8824 2146 8895
rect 2272 8824 2304 8895
rect 2430 8824 2462 8895
rect 2588 8824 2620 8895
rect 2746 8824 2778 8895
rect 2904 8824 2936 8895
rect 3062 8824 3094 8895
rect 3220 8824 3252 8895
rect 3378 8824 3410 8895
rect 3536 8824 3568 8895
rect 3694 8824 3726 8895
rect 505 8787 3765 8824
rect 505 8782 671 8787
rect 505 8500 552 8782
rect 505 8496 671 8500
rect 692 8496 724 8787
rect 850 8496 882 8787
rect 1008 8496 1040 8787
rect 1166 8496 1198 8787
rect 1324 8496 1356 8787
rect 1482 8496 1514 8787
rect 1640 8496 1672 8787
rect 1798 8496 1830 8787
rect 1956 8496 1988 8787
rect 2114 8496 2146 8787
rect 2272 8496 2304 8787
rect 2430 8496 2462 8787
rect 2588 8496 2620 8787
rect 2746 8496 2778 8787
rect 2904 8496 2936 8787
rect 3062 8496 3094 8787
rect 3220 8496 3252 8787
rect 3378 8496 3410 8787
rect 3536 8496 3568 8787
rect 3694 8496 3726 8787
rect 505 8459 3757 8496
rect 505 8454 671 8459
rect 505 8392 552 8454
rect 505 8388 671 8392
rect 692 8388 724 8459
rect 850 8388 882 8459
rect 1008 8388 1040 8459
rect 1166 8388 1198 8459
rect 1324 8388 1356 8459
rect 1482 8388 1514 8459
rect 1640 8388 1672 8459
rect 1798 8388 1830 8459
rect 1956 8388 1988 8459
rect 2114 8388 2146 8459
rect 2272 8388 2304 8459
rect 2430 8388 2462 8459
rect 2588 8388 2620 8459
rect 2746 8388 2778 8459
rect 2904 8388 2936 8459
rect 3062 8388 3094 8459
rect 3220 8388 3252 8459
rect 3378 8388 3410 8459
rect 3536 8388 3568 8459
rect 3694 8388 3726 8459
rect 505 8351 3765 8388
rect 505 8346 671 8351
rect 505 8064 552 8346
rect 505 8060 671 8064
rect 692 8060 724 8351
rect 850 8060 882 8351
rect 1008 8060 1040 8351
rect 1166 8060 1198 8351
rect 1324 8060 1356 8351
rect 1482 8060 1514 8351
rect 1640 8060 1672 8351
rect 1798 8060 1830 8351
rect 1956 8060 1988 8351
rect 2114 8060 2146 8351
rect 2272 8060 2304 8351
rect 2430 8060 2462 8351
rect 2588 8060 2620 8351
rect 2746 8060 2778 8351
rect 2904 8060 2936 8351
rect 3062 8060 3094 8351
rect 3220 8060 3252 8351
rect 3378 8060 3410 8351
rect 3536 8060 3568 8351
rect 3694 8060 3726 8351
rect 505 8023 3757 8060
rect 505 8018 671 8023
rect 505 7956 552 8018
rect 505 7952 671 7956
rect 692 7952 724 8023
rect 850 7952 882 8023
rect 1008 7952 1040 8023
rect 1166 7952 1198 8023
rect 1324 7952 1356 8023
rect 1482 7952 1514 8023
rect 1640 7952 1672 8023
rect 1798 7952 1830 8023
rect 1956 7952 1988 8023
rect 2114 7952 2146 8023
rect 2272 7952 2304 8023
rect 2430 7952 2462 8023
rect 2588 7952 2620 8023
rect 2746 7952 2778 8023
rect 2904 7952 2936 8023
rect 3062 7952 3094 8023
rect 3220 7952 3252 8023
rect 3378 7952 3410 8023
rect 3536 7952 3568 8023
rect 3694 7952 3726 8023
rect 505 7915 3765 7952
rect 505 7910 671 7915
rect 505 7628 552 7910
rect 505 7624 671 7628
rect 692 7624 724 7915
rect 850 7624 882 7915
rect 1008 7624 1040 7915
rect 1166 7624 1198 7915
rect 1324 7624 1356 7915
rect 1482 7624 1514 7915
rect 1640 7624 1672 7915
rect 1798 7624 1830 7915
rect 1956 7624 1988 7915
rect 2114 7624 2146 7915
rect 2272 7624 2304 7915
rect 2430 7624 2462 7915
rect 2588 7624 2620 7915
rect 2746 7624 2778 7915
rect 2904 7624 2936 7915
rect 3062 7624 3094 7915
rect 3220 7624 3252 7915
rect 3378 7624 3410 7915
rect 3536 7624 3568 7915
rect 3694 7624 3726 7915
rect 505 7587 3757 7624
rect 505 7582 671 7587
rect 505 7520 552 7582
rect 505 7516 671 7520
rect 692 7516 724 7587
rect 850 7516 882 7587
rect 1008 7516 1040 7587
rect 1166 7516 1198 7587
rect 1324 7516 1356 7587
rect 1482 7516 1514 7587
rect 1640 7516 1672 7587
rect 1798 7516 1830 7587
rect 1956 7516 1988 7587
rect 2114 7516 2146 7587
rect 2272 7516 2304 7587
rect 2430 7516 2462 7587
rect 2588 7516 2620 7587
rect 2746 7516 2778 7587
rect 2904 7516 2936 7587
rect 3062 7516 3094 7587
rect 3220 7516 3252 7587
rect 3378 7516 3410 7587
rect 3536 7516 3568 7587
rect 3694 7516 3726 7587
rect 505 7479 3765 7516
rect 505 7474 671 7479
rect 505 7192 552 7474
rect 505 7188 671 7192
rect 692 7188 724 7479
rect 850 7188 882 7479
rect 1008 7188 1040 7479
rect 1166 7188 1198 7479
rect 1324 7188 1356 7479
rect 1482 7188 1514 7479
rect 1640 7188 1672 7479
rect 1798 7188 1830 7479
rect 1956 7188 1988 7479
rect 2114 7188 2146 7479
rect 2272 7188 2304 7479
rect 2430 7188 2462 7479
rect 2588 7188 2620 7479
rect 2746 7188 2778 7479
rect 2904 7188 2936 7479
rect 3062 7188 3094 7479
rect 3220 7188 3252 7479
rect 3378 7188 3410 7479
rect 3536 7188 3568 7479
rect 3694 7188 3726 7479
rect 505 7151 3757 7188
rect 505 7146 671 7151
rect 505 7084 552 7146
rect 505 7080 671 7084
rect 692 7080 724 7151
rect 850 7080 882 7151
rect 1008 7080 1040 7151
rect 1166 7080 1198 7151
rect 1324 7080 1356 7151
rect 1482 7080 1514 7151
rect 1640 7080 1672 7151
rect 1798 7080 1830 7151
rect 1956 7080 1988 7151
rect 2114 7080 2146 7151
rect 2272 7080 2304 7151
rect 2430 7080 2462 7151
rect 2588 7080 2620 7151
rect 2746 7080 2778 7151
rect 2904 7080 2936 7151
rect 3062 7080 3094 7151
rect 3220 7080 3252 7151
rect 3378 7080 3410 7151
rect 3536 7080 3568 7151
rect 3694 7080 3726 7151
rect 505 7043 3765 7080
rect 505 7038 671 7043
rect 505 6756 552 7038
rect 505 6752 671 6756
rect 692 6752 724 7043
rect 850 6752 882 7043
rect 1008 6752 1040 7043
rect 1166 6752 1198 7043
rect 1324 6752 1356 7043
rect 1482 6752 1514 7043
rect 1640 6752 1672 7043
rect 1798 6752 1830 7043
rect 1956 6752 1988 7043
rect 2114 6752 2146 7043
rect 2272 6752 2304 7043
rect 2430 6752 2462 7043
rect 2588 6752 2620 7043
rect 2746 6752 2778 7043
rect 2904 6752 2936 7043
rect 3062 6752 3094 7043
rect 3220 6752 3252 7043
rect 3378 6752 3410 7043
rect 3536 6752 3568 7043
rect 3694 6752 3726 7043
rect 505 6715 3757 6752
rect 505 6710 671 6715
rect 505 6648 552 6710
rect 505 6644 671 6648
rect 692 6644 724 6715
rect 850 6644 882 6715
rect 1008 6644 1040 6715
rect 1166 6644 1198 6715
rect 1324 6644 1356 6715
rect 1482 6644 1514 6715
rect 1640 6644 1672 6715
rect 1798 6644 1830 6715
rect 1956 6644 1988 6715
rect 2114 6644 2146 6715
rect 2272 6644 2304 6715
rect 2430 6644 2462 6715
rect 2588 6644 2620 6715
rect 2746 6644 2778 6715
rect 2904 6644 2936 6715
rect 3062 6644 3094 6715
rect 3220 6644 3252 6715
rect 3378 6644 3410 6715
rect 3536 6644 3568 6715
rect 3694 6644 3726 6715
rect 505 6607 3765 6644
rect 505 6602 671 6607
rect 505 6320 552 6602
rect 505 6316 671 6320
rect 692 6316 724 6607
rect 850 6316 882 6607
rect 1008 6316 1040 6607
rect 1166 6316 1198 6607
rect 1324 6316 1356 6607
rect 1482 6316 1514 6607
rect 1640 6316 1672 6607
rect 1798 6316 1830 6607
rect 1956 6316 1988 6607
rect 2114 6316 2146 6607
rect 2272 6316 2304 6607
rect 2430 6316 2462 6607
rect 2588 6316 2620 6607
rect 2746 6316 2778 6607
rect 2904 6316 2936 6607
rect 3062 6316 3094 6607
rect 3220 6316 3252 6607
rect 3378 6316 3410 6607
rect 3536 6316 3568 6607
rect 3694 6316 3726 6607
rect 505 6279 3757 6316
rect 505 6274 671 6279
rect 505 6212 552 6274
rect 505 6208 671 6212
rect 692 6208 724 6279
rect 850 6208 882 6279
rect 1008 6208 1040 6279
rect 1166 6208 1198 6279
rect 1324 6208 1356 6279
rect 1482 6208 1514 6279
rect 1640 6208 1672 6279
rect 1798 6208 1830 6279
rect 1956 6208 1988 6279
rect 2114 6208 2146 6279
rect 2272 6208 2304 6279
rect 2430 6208 2462 6279
rect 2588 6208 2620 6279
rect 2746 6208 2778 6279
rect 2904 6208 2936 6279
rect 3062 6208 3094 6279
rect 3220 6208 3252 6279
rect 3378 6208 3410 6279
rect 3536 6208 3568 6279
rect 3694 6208 3726 6279
rect 505 6171 3765 6208
rect 505 6166 671 6171
rect 505 5884 552 6166
rect 505 5880 671 5884
rect 692 5880 724 6171
rect 850 5880 882 6171
rect 1008 5880 1040 6171
rect 1166 5880 1198 6171
rect 1324 5880 1356 6171
rect 1482 5880 1514 6171
rect 1640 5880 1672 6171
rect 1798 5880 1830 6171
rect 1956 5880 1988 6171
rect 2114 5880 2146 6171
rect 2272 5880 2304 6171
rect 2430 5880 2462 6171
rect 2588 5880 2620 6171
rect 2746 5880 2778 6171
rect 2904 5880 2936 6171
rect 3062 5880 3094 6171
rect 3220 5880 3252 6171
rect 3378 5880 3410 6171
rect 3536 5880 3568 6171
rect 3694 5880 3726 6171
rect 505 5843 3757 5880
rect 505 5838 671 5843
rect 505 5776 552 5838
rect 505 5772 671 5776
rect 692 5772 724 5843
rect 850 5772 882 5843
rect 1008 5772 1040 5843
rect 1166 5772 1198 5843
rect 1324 5772 1356 5843
rect 1482 5772 1514 5843
rect 1640 5772 1672 5843
rect 1798 5772 1830 5843
rect 1956 5772 1988 5843
rect 2114 5772 2146 5843
rect 2272 5772 2304 5843
rect 2430 5772 2462 5843
rect 2588 5772 2620 5843
rect 2746 5772 2778 5843
rect 2904 5772 2936 5843
rect 3062 5772 3094 5843
rect 3220 5772 3252 5843
rect 3378 5772 3410 5843
rect 3536 5772 3568 5843
rect 3694 5772 3726 5843
rect 505 5735 3765 5772
rect 505 5730 671 5735
rect 505 5448 552 5730
rect 505 5444 671 5448
rect 692 5444 724 5735
rect 850 5444 882 5735
rect 1008 5444 1040 5735
rect 1166 5444 1198 5735
rect 1324 5444 1356 5735
rect 1482 5444 1514 5735
rect 1640 5444 1672 5735
rect 1798 5444 1830 5735
rect 1956 5444 1988 5735
rect 2114 5444 2146 5735
rect 2272 5444 2304 5735
rect 2430 5444 2462 5735
rect 2588 5444 2620 5735
rect 2746 5444 2778 5735
rect 2904 5444 2936 5735
rect 3062 5444 3094 5735
rect 3220 5444 3252 5735
rect 3378 5444 3410 5735
rect 3536 5444 3568 5735
rect 3694 5444 3726 5735
rect 505 5407 3757 5444
rect 505 5402 671 5407
rect 505 5340 552 5402
rect 505 5336 671 5340
rect 692 5336 724 5407
rect 850 5336 882 5407
rect 1008 5336 1040 5407
rect 1166 5336 1198 5407
rect 1324 5336 1356 5407
rect 1482 5336 1514 5407
rect 1640 5336 1672 5407
rect 1798 5336 1830 5407
rect 1956 5336 1988 5407
rect 2114 5336 2146 5407
rect 2272 5336 2304 5407
rect 2430 5336 2462 5407
rect 2588 5336 2620 5407
rect 2746 5336 2778 5407
rect 2904 5336 2936 5407
rect 3062 5336 3094 5407
rect 3220 5336 3252 5407
rect 3378 5336 3410 5407
rect 3536 5336 3568 5407
rect 3694 5336 3726 5407
rect 505 5299 3765 5336
rect 505 5294 671 5299
rect 505 5012 552 5294
rect 505 5008 671 5012
rect 692 5008 724 5299
rect 850 5008 882 5299
rect 1008 5008 1040 5299
rect 1166 5008 1198 5299
rect 1324 5008 1356 5299
rect 1482 5008 1514 5299
rect 1640 5008 1672 5299
rect 1798 5008 1830 5299
rect 1956 5008 1988 5299
rect 2114 5008 2146 5299
rect 2272 5008 2304 5299
rect 2430 5008 2462 5299
rect 2588 5008 2620 5299
rect 2746 5008 2778 5299
rect 2904 5008 2936 5299
rect 3062 5008 3094 5299
rect 3220 5008 3252 5299
rect 3378 5008 3410 5299
rect 3536 5008 3568 5299
rect 3694 5008 3726 5299
rect 505 4971 3757 5008
rect 505 4966 671 4971
rect 505 4904 552 4966
rect 505 4900 671 4904
rect 692 4900 724 4971
rect 850 4900 882 4971
rect 1008 4900 1040 4971
rect 1166 4900 1198 4971
rect 1324 4900 1356 4971
rect 1482 4900 1514 4971
rect 1640 4900 1672 4971
rect 1798 4900 1830 4971
rect 1956 4900 1988 4971
rect 2114 4900 2146 4971
rect 2272 4900 2304 4971
rect 2430 4900 2462 4971
rect 2588 4900 2620 4971
rect 2746 4900 2778 4971
rect 2904 4900 2936 4971
rect 3062 4900 3094 4971
rect 3220 4900 3252 4971
rect 3378 4900 3410 4971
rect 3536 4900 3568 4971
rect 3694 4900 3726 4971
rect 505 4863 3765 4900
rect 505 4858 671 4863
rect 505 4576 552 4858
rect 505 4572 671 4576
rect 692 4572 724 4863
rect 850 4572 882 4863
rect 1008 4572 1040 4863
rect 1166 4572 1198 4863
rect 1324 4572 1356 4863
rect 1482 4572 1514 4863
rect 1640 4572 1672 4863
rect 1798 4572 1830 4863
rect 1956 4572 1988 4863
rect 2114 4572 2146 4863
rect 2272 4572 2304 4863
rect 2430 4572 2462 4863
rect 2588 4572 2620 4863
rect 2746 4572 2778 4863
rect 2904 4572 2936 4863
rect 3062 4572 3094 4863
rect 3220 4572 3252 4863
rect 3378 4572 3410 4863
rect 3536 4572 3568 4863
rect 3694 4572 3726 4863
rect 505 4535 3755 4572
rect 505 4530 671 4535
rect 850 4530 882 4535
rect 1008 4530 1040 4535
rect 1166 4530 1198 4535
rect 1324 4530 1356 4535
rect 1482 4530 1514 4535
rect 1640 4530 1672 4535
rect 1798 4530 1830 4535
rect 1956 4530 1988 4535
rect 2114 4530 2146 4535
rect 2272 4530 2304 4535
rect 2430 4530 2462 4535
rect 2588 4530 2620 4535
rect 2746 4530 2778 4535
rect 2904 4530 2936 4535
rect 3062 4530 3094 4535
rect 3220 4530 3252 4535
rect 3378 4530 3410 4535
rect 3536 4530 3568 4535
rect 3694 4530 3726 4535
rect 505 3756 552 4530
rect 599 4452 3820 4472
rect 599 4390 639 4452
rect 3787 4440 3820 4452
rect 3790 4398 3820 4440
rect 3787 4390 3820 4398
rect 599 4373 3820 4390
rect 692 4294 724 4300
rect 850 4294 882 4300
rect 1008 4294 1040 4300
rect 1166 4294 1198 4300
rect 1324 4294 1356 4300
rect 1482 4294 1514 4300
rect 1640 4294 1672 4300
rect 1798 4294 1830 4300
rect 1956 4294 1988 4300
rect 2114 4294 2146 4300
rect 2272 4294 2304 4300
rect 2430 4294 2462 4300
rect 2588 4294 2620 4300
rect 2746 4294 2778 4300
rect 2904 4294 2936 4300
rect 3062 4294 3094 4300
rect 3220 4294 3252 4300
rect 3378 4294 3410 4300
rect 3536 4294 3568 4300
rect 3694 4294 3726 4300
rect 654 4257 3765 4294
rect 692 3967 724 4257
rect 850 3967 882 4257
rect 1008 3967 1040 4257
rect 1166 3967 1198 4257
rect 1324 3967 1356 4257
rect 1482 3967 1514 4257
rect 1640 3967 1672 4257
rect 1798 3967 1830 4257
rect 1956 3967 1988 4257
rect 2114 3967 2146 4257
rect 2272 3967 2304 4257
rect 2430 3967 2462 4257
rect 2588 3967 2620 4257
rect 2746 3967 2778 4257
rect 2904 3967 2936 4257
rect 3062 3967 3094 4257
rect 3220 3967 3252 4257
rect 3378 3967 3410 4257
rect 3536 3967 3568 4257
rect 3694 3967 3726 4257
rect 651 3930 3762 3967
rect 692 3926 724 3930
rect 850 3926 882 3930
rect 1008 3926 1040 3930
rect 1166 3926 1198 3930
rect 1324 3926 1356 3930
rect 1482 3926 1514 3930
rect 1640 3926 1672 3930
rect 1798 3926 1830 3930
rect 1956 3926 1988 3930
rect 2114 3926 2146 3930
rect 2272 3926 2304 3930
rect 2430 3926 2462 3930
rect 2588 3926 2620 3930
rect 2746 3926 2778 3930
rect 2904 3926 2936 3930
rect 651 3841 2959 3856
rect 651 3806 677 3841
rect 2924 3806 2959 3841
rect 651 3792 2959 3806
rect 505 3709 2158 3756
rect 446 3665 2040 3671
rect 446 3617 475 3665
rect 2008 3617 2040 3665
rect 446 3610 2040 3617
rect 446 3385 457 3610
rect 2111 3540 2158 3709
rect 2203 3666 2980 3673
rect 2203 3619 2232 3666
rect 2946 3619 2980 3666
rect 2203 3605 2980 3619
rect 3015 3540 3053 3930
rect 3062 3926 3094 3930
rect 3220 3926 3252 3930
rect 3378 3926 3410 3930
rect 3536 3926 3568 3930
rect 3694 3926 3726 3930
rect 3910 3855 3930 10644
rect 3093 3839 3930 3855
rect 3093 3805 3114 3839
rect 3806 3805 3930 3839
rect 3093 3792 3930 3805
rect 3910 3672 3930 3792
rect 3096 3662 3930 3672
rect 3096 3615 3123 3662
rect 3799 3615 3930 3662
rect 3096 3605 3930 3615
rect 2091 3521 2179 3540
rect 350 1183 457 3385
rect 591 3188 628 3435
rect 687 3188 718 3497
rect 845 3188 876 3497
rect 1003 3188 1034 3497
rect 591 3150 1074 3188
rect 502 1401 549 2628
rect 587 1831 627 2724
rect 686 2090 723 3150
rect 1429 3097 1460 3499
rect 1587 3097 1618 3508
rect 866 3066 1618 3097
rect 1587 2908 1618 3066
rect 1745 2974 1776 3512
rect 1903 2974 1934 3512
rect 2091 3105 2107 3521
rect 2166 3105 2179 3521
rect 2995 3524 3072 3540
rect 2329 3191 2360 3498
rect 2487 3191 2518 3498
rect 2645 3191 2676 3498
rect 2714 3191 2765 3234
rect 2803 3191 2834 3498
rect 2295 3148 2873 3191
rect 2091 3089 2179 3105
rect 2995 3101 3006 3524
rect 3061 3101 3072 3524
rect 3231 3189 3262 3504
rect 3389 3189 3420 3504
rect 3547 3191 3578 3504
rect 3618 3191 3664 3266
rect 3705 3191 3736 3504
rect 3516 3189 3766 3191
rect 3198 3148 3770 3189
rect 3516 3145 3766 3148
rect 3910 3128 3930 3605
rect 3969 4498 4014 10703
rect 4087 4498 4124 10827
rect 3969 4380 4124 4498
rect 3969 3697 4014 4380
rect 4087 3697 4124 4380
rect 3969 3588 4124 3697
rect 3969 3128 4014 3588
rect 3910 3102 4014 3128
rect 2995 3087 3072 3101
rect 4087 3082 4124 3588
rect 4167 3082 4188 10827
rect 4087 3055 4188 3082
rect 3919 2991 4153 2999
rect 3000 2974 3031 2975
rect 3919 2974 3928 2991
rect 1745 2943 3928 2974
rect 1587 2877 2794 2908
rect 811 2659 969 2661
rect 811 2615 1398 2659
rect 811 2614 969 2615
rect 846 2613 969 2614
rect 1246 2613 1398 2615
rect 846 2312 877 2613
rect 1276 2310 1307 2613
rect 1346 2586 1398 2613
rect 1705 2311 1736 2877
rect 1863 2794 2178 2825
rect 1863 2345 1894 2794
rect 2294 2639 2325 2653
rect 1846 2308 1909 2345
rect 821 2221 2256 2242
rect 821 2170 864 2221
rect 2214 2170 2256 2221
rect 821 2151 2256 2170
rect 2293 2200 2328 2639
rect 2763 2314 2794 2877
rect 3000 2652 3031 2943
rect 3919 2925 3928 2943
rect 4143 2925 4153 2991
rect 3919 2917 4153 2925
rect 3784 2804 4157 2831
rect 3000 2313 3034 2652
rect 3000 2309 3031 2313
rect 3473 2200 3504 2651
rect 3631 2200 3662 2651
rect 2293 2165 3662 2200
rect 3784 2196 3824 2804
rect 3879 2196 4157 2804
rect 686 2053 2868 2090
rect 678 2004 2773 2017
rect 678 1952 725 2004
rect 2739 2000 2773 2004
rect 2742 1963 2773 2000
rect 2739 1952 2773 1963
rect 678 1923 2773 1952
rect 678 1916 935 1923
rect 587 1791 805 1831
rect 752 1281 788 1567
rect 893 1508 935 1916
rect 892 1443 935 1508
rect 973 1916 2773 1923
rect 973 1910 1193 1916
rect 973 1443 1110 1910
rect 892 1442 1110 1443
rect 1151 1449 1193 1910
rect 1362 1817 1928 1863
rect 1464 1785 1510 1817
rect 1780 1785 1826 1817
rect 1391 1553 1422 1776
rect 1549 1553 1580 1776
rect 1707 1553 1738 1776
rect 1865 1553 1896 1776
rect 1151 1442 2240 1449
rect 892 1419 2240 1442
rect 892 1371 1297 1419
rect 2190 1371 2240 1419
rect 892 1336 2240 1371
rect 892 1203 1193 1336
rect 2295 1281 2326 1855
rect 2399 1307 2462 1780
rect 2526 1385 2654 1786
rect 2725 1516 2756 1825
rect 2831 1584 2868 2053
rect 2940 1625 2975 2165
rect 3784 2094 4157 2196
rect 3093 2077 4157 2094
rect 3093 1938 3121 2077
rect 3813 1987 4157 2077
rect 3813 1938 3825 1987
rect 3093 1914 3825 1938
rect 3154 1440 3185 1856
rect 3312 1440 3343 1856
rect 3470 1440 3501 1856
rect 3628 1539 3659 1856
rect 3627 1517 3659 1539
rect 3627 1440 3658 1517
rect 3154 1434 3658 1440
rect 3154 1409 3169 1434
rect 3155 1382 3169 1409
rect 3634 1409 3658 1434
rect 3634 1382 3643 1409
rect 3155 1372 3643 1382
rect 3784 1379 3825 1914
rect 3880 1379 4157 1987
rect 3784 1338 4157 1379
rect 2399 1244 3764 1307
rect 350 886 360 1183
rect 447 886 457 1183
rect 509 1180 3369 1203
rect 509 1117 553 1180
rect 3320 1117 3369 1180
rect 509 1095 3369 1117
rect 350 864 457 886
rect 430 742 537 779
rect 604 772 1036 1008
rect 3437 964 3764 1244
rect 3943 1204 4157 1338
rect 3943 1183 4004 1204
rect 430 597 459 742
rect 506 597 537 742
rect 430 548 537 597
rect 588 667 1024 682
rect 588 612 605 667
rect 1008 612 1024 667
rect 588 596 1024 612
rect 3337 606 3769 842
rect 3943 548 3960 1183
rect 383 524 3960 548
rect 383 463 406 524
rect 3940 519 3960 524
rect 4000 519 4004 1183
rect 3940 508 4004 519
rect 4058 508 4157 1204
rect 3940 463 4157 508
rect 383 442 4157 463
rect 179 281 283 292
rect 179 253 4195 281
rect 179 199 255 253
rect 4117 199 4195 253
rect 179 169 4195 199
rect 4278 102 4301 11029
rect 0 72 4301 102
rect 0 26 148 72
rect 4259 70 4301 72
rect 4347 70 4377 11078
rect 4259 26 4377 70
rect 0 0 4377 26
<< via1 >>
rect 544 10706 3758 10718
rect 544 10671 3758 10706
rect 544 10664 3758 10671
rect 360 10410 446 10428
rect 360 3817 383 10410
rect 383 3817 437 10410
rect 437 3817 446 10410
rect 360 3385 446 3817
rect 639 4440 3787 4452
rect 639 4398 646 4440
rect 646 4398 3787 4440
rect 639 4390 3787 4398
rect 2107 3105 2166 3521
rect 3006 3101 3061 3524
rect 3928 2925 4143 2991
rect 725 2000 2739 2004
rect 725 1963 734 2000
rect 734 1963 2739 2000
rect 725 1952 2739 1963
rect 3121 1938 3813 2077
rect 3169 1382 3634 1434
rect 360 886 447 1183
rect 553 1169 3320 1180
rect 553 1133 564 1169
rect 564 1133 3290 1169
rect 3290 1133 3320 1169
rect 553 1117 3320 1133
rect 605 612 1008 667
rect 406 516 3940 524
rect 406 479 454 516
rect 454 479 3919 516
rect 3919 479 3940 516
rect 4004 508 4058 1204
rect 406 463 3940 479
<< metal2 >>
rect 257 10718 3800 10782
rect 257 10664 544 10718
rect 3758 10664 3800 10718
rect 257 10624 3800 10664
rect 257 10428 549 10624
rect 3861 10579 4153 10782
rect 596 10450 4153 10579
rect 257 3605 360 10428
rect 258 3385 360 3605
rect 446 10320 549 10428
rect 446 10191 3825 10320
rect 446 9884 549 10191
rect 3861 10143 4153 10450
rect 596 10014 4153 10143
rect 446 9755 3825 9884
rect 446 9448 549 9755
rect 3861 9707 4153 10014
rect 596 9578 4153 9707
rect 446 9319 3825 9448
rect 446 9012 549 9319
rect 3861 9271 4153 9578
rect 596 9142 4153 9271
rect 446 8883 3825 9012
rect 446 8576 549 8883
rect 3861 8835 4153 9142
rect 596 8706 4153 8835
rect 446 8447 3825 8576
rect 446 8140 549 8447
rect 3861 8399 4153 8706
rect 596 8270 4153 8399
rect 446 8011 3825 8140
rect 446 7704 549 8011
rect 3861 7963 4153 8270
rect 596 7834 4153 7963
rect 446 7575 3825 7704
rect 446 7268 549 7575
rect 3861 7527 4153 7834
rect 596 7398 4153 7527
rect 446 7139 3825 7268
rect 446 6832 549 7139
rect 3861 7091 4153 7398
rect 596 6962 4153 7091
rect 446 6703 3825 6832
rect 446 6396 549 6703
rect 3861 6655 4153 6962
rect 596 6526 4153 6655
rect 446 6267 3825 6396
rect 446 5960 549 6267
rect 3861 6219 4153 6526
rect 596 6090 4153 6219
rect 446 5831 3825 5960
rect 446 5524 549 5831
rect 3861 5783 4153 6090
rect 596 5654 4153 5783
rect 446 5395 3825 5524
rect 446 5088 549 5395
rect 3861 5347 4153 5654
rect 596 5218 4153 5347
rect 446 4959 3825 5088
rect 446 4652 549 4959
rect 3861 4911 4153 5218
rect 596 4782 4153 4911
rect 446 4523 3825 4652
rect 446 4475 549 4523
rect 446 4452 3823 4475
rect 446 4390 639 4452
rect 3787 4390 3823 4452
rect 446 4369 3823 4390
rect 446 4048 549 4369
rect 3861 4307 4153 4782
rect 599 4178 4153 4307
rect 446 3919 3828 4048
rect 446 3855 549 3919
rect 3861 3875 4153 4178
rect 446 3778 3829 3855
rect 446 3605 3828 3778
rect 446 3463 549 3605
rect 2091 3521 2179 3540
rect 446 3462 558 3463
rect 446 3385 1148 3462
rect 258 3375 1148 3385
rect 1205 3376 2043 3460
rect 1205 3289 1289 3376
rect 573 3205 1289 3289
rect 257 3110 457 3180
rect 1493 3112 1556 3348
rect 257 3048 864 3110
rect 1101 3049 1556 3112
rect 257 2980 457 3048
rect 583 2836 626 3048
rect 1101 2860 1164 3049
rect 1802 2987 1865 3348
rect 2091 3109 2107 3521
rect 910 2797 1164 2860
rect 1340 2924 1865 2987
rect 2004 3105 2107 3109
rect 2166 3109 2179 3521
rect 2210 3462 2295 3605
rect 2995 3524 3072 3540
rect 2210 3377 2934 3462
rect 2392 3109 2458 3348
rect 2166 3105 2458 3109
rect 2004 3043 2458 3105
rect 910 2661 973 2797
rect 526 2596 973 2661
rect 729 2259 841 2526
rect 910 2460 973 2596
rect 1151 2259 1263 2527
rect 1340 2458 1403 2924
rect 2004 2876 2070 3043
rect 2707 2956 2773 3349
rect 2995 3107 3006 3524
rect 1609 2810 2070 2876
rect 2159 2828 2213 2956
rect 2322 2890 2773 2956
rect 2912 3101 3006 3107
rect 3061 3107 3072 3524
rect 3110 3462 3195 3605
rect 3110 3377 3834 3462
rect 3110 3376 3197 3377
rect 3133 3317 3139 3376
rect 3191 3317 3197 3376
rect 3292 3107 3358 3348
rect 3449 3317 3455 3377
rect 3507 3317 3513 3377
rect 3061 3101 3358 3107
rect 2912 3041 3358 3101
rect 1609 2456 1675 2810
rect 2322 2742 2388 2890
rect 1930 2676 2388 2742
rect 1742 2413 1854 2526
rect 1930 2454 1996 2676
rect 2912 2632 2978 3041
rect 3607 2947 3673 3349
rect 3766 3317 3772 3377
rect 3824 3317 3830 3377
rect 2621 2566 2978 2632
rect 3105 2881 3673 2947
rect 3919 2991 4153 3875
rect 3919 2925 3928 2991
rect 4143 2925 4153 2991
rect 1742 2323 2264 2413
rect 2343 2259 2446 2514
rect 2621 2462 2687 2566
rect 2845 2413 2957 2527
rect 3105 2460 3171 2881
rect 3238 2557 3748 2647
rect 3238 2413 3328 2557
rect 2845 2323 3328 2413
rect 3514 2259 3617 2513
rect 259 2077 3832 2259
rect 259 2004 3121 2077
rect 259 1952 725 2004
rect 2739 1952 3121 2004
rect 259 1938 3121 1952
rect 3813 1938 3832 2077
rect 259 1741 3832 1938
rect 3919 1623 4153 2925
rect 1228 1510 3000 1623
rect 3078 1510 4153 1623
rect 261 1283 461 1447
rect 551 1434 3649 1445
rect 551 1401 3169 1434
rect 3148 1382 3169 1401
rect 3634 1401 3649 1434
rect 3634 1382 3648 1401
rect 3148 1381 3648 1382
rect 261 1247 2326 1283
rect 3943 1204 4157 1284
rect 3943 1203 4004 1204
rect 350 1183 457 1203
rect 350 886 360 1183
rect 447 886 457 1183
rect 509 1180 4004 1203
rect 509 1117 553 1180
rect 3320 1117 4004 1180
rect 509 1095 4004 1117
rect 350 682 457 886
rect 350 667 1024 682
rect 350 612 605 667
rect 1008 612 1024 667
rect 350 598 1024 612
rect 3943 548 4004 1095
rect 383 524 4004 548
rect 383 463 406 524
rect 3940 508 4004 524
rect 4058 508 4157 1204
rect 3940 463 4157 508
rect 383 442 4157 463
use amp_via_2cut  amp_via_2cut_0
timestamp 1717613630
transform 0 1 8530 -1 0 20917
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_1
timestamp 1717613630
transform 0 1 8688 -1 0 20829
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_2
timestamp 1717613630
transform 0 1 9004 -1 0 20829
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_3
timestamp 1717613630
transform 0 1 8846 -1 0 20917
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_4
timestamp 1717613630
transform 0 1 10584 -1 0 20224
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_5
timestamp 1717613630
transform 0 1 10426 -1 0 20312
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_6
timestamp 1717613630
transform 0 1 9320 -1 0 20224
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_7
timestamp 1717613630
transform 0 1 9162 -1 0 20312
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_8
timestamp 1717613630
transform 0 1 9636 -1 0 20224
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_9
timestamp 1717613630
transform 0 1 9478 -1 0 20312
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_10
timestamp 1717613630
transform 0 1 9952 -1 0 20224
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_11
timestamp 1717613630
transform 0 1 9794 -1 0 20312
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_12
timestamp 1717613630
transform 0 1 10268 -1 0 20224
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_13
timestamp 1717613630
transform 0 1 10110 -1 0 20312
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_14
timestamp 1717613630
transform 0 1 11532 -1 0 20829
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_15
timestamp 1717613630
transform 0 1 11690 -1 0 20917
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_16
timestamp 1717613630
transform 0 1 10900 -1 0 20829
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_17
timestamp 1717613630
transform 0 1 10742 -1 0 20917
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_18
timestamp 1717613630
transform 0 1 11216 -1 0 20829
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_19
timestamp 1717613630
transform 0 1 11058 -1 0 20917
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_20
timestamp 1717613630
transform 0 1 11374 -1 0 20917
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_21
timestamp 1717613630
transform 0 1 9004 -1 0 20224
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_22
timestamp 1717613630
transform 0 1 8846 -1 0 20312
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_23
timestamp 1717613630
transform 0 1 8530 -1 0 20312
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_24
timestamp 1717613630
transform 0 1 8999 1 0 -12777
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_25
timestamp 1717613630
transform 0 1 9478 -1 0 20917
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_26
timestamp 1717613630
transform 0 1 9162 -1 0 20917
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_27
timestamp 1717613630
transform 0 1 9320 -1 0 20829
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_28
timestamp 1717613630
transform 0 1 9794 -1 0 20917
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_29
timestamp 1717613630
transform 0 1 9952 -1 0 20829
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_30
timestamp 1717613630
transform 0 1 9636 -1 0 20829
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_31
timestamp 1717613630
transform 0 1 10426 -1 0 20917
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_32
timestamp 1717613630
transform 0 1 10268 -1 0 20829
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_33
timestamp 1717613630
transform 0 1 10110 -1 0 20917
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_34
timestamp 1717613630
transform 0 1 10584 -1 0 20829
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_35
timestamp 1717613630
transform 0 1 11690 -1 0 20312
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_36
timestamp 1717613630
transform 0 1 11532 -1 0 20224
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_37
timestamp 1717613630
transform 0 1 11374 -1 0 20312
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_38
timestamp 1717613630
transform 0 1 11216 -1 0 20224
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_39
timestamp 1717613630
transform 0 1 11058 -1 0 20312
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_40
timestamp 1717613630
transform 0 1 10900 -1 0 20224
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_41
timestamp 1717613630
transform 0 1 10742 -1 0 20312
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_42
timestamp 1717613630
transform 0 1 8846 -1 0 21353
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_43
timestamp 1717613630
transform 0 1 9004 -1 0 21265
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_44
timestamp 1717613630
transform 0 1 8530 -1 0 21353
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_45
timestamp 1717613630
transform 0 1 8688 -1 0 21265
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_46
timestamp 1717613630
transform 0 1 10584 -1 0 21265
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_47
timestamp 1717613630
transform 0 1 10426 -1 0 21353
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_48
timestamp 1717613630
transform 0 1 10268 -1 0 21265
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_49
timestamp 1717613630
transform 0 1 10110 -1 0 21353
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_50
timestamp 1717613630
transform 0 1 9794 -1 0 21353
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_51
timestamp 1717613630
transform 0 1 9952 -1 0 21265
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_52
timestamp 1717613630
transform 0 1 9478 -1 0 21353
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_53
timestamp 1717613630
transform 0 1 9636 -1 0 21265
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_54
timestamp 1717613630
transform 0 1 9162 -1 0 21353
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_55
timestamp 1717613630
transform 0 1 9320 -1 0 21265
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_56
timestamp 1717613630
transform 0 1 11690 -1 0 21353
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_57
timestamp 1717613630
transform 0 1 11532 -1 0 21265
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_58
timestamp 1717613630
transform 0 1 11374 -1 0 21353
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_59
timestamp 1717613630
transform 0 1 11216 -1 0 21265
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_60
timestamp 1717613630
transform 0 1 11058 -1 0 21353
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_61
timestamp 1717613630
transform 0 1 10900 -1 0 21265
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_62
timestamp 1717613630
transform 0 1 10742 -1 0 21353
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_63
timestamp 1717613630
transform 0 1 11690 -1 0 22661
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_64
timestamp 1717613630
transform 0 1 11532 -1 0 22573
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_65
timestamp 1717613630
transform 0 1 11374 -1 0 22661
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_66
timestamp 1717613630
transform 0 1 11216 -1 0 22573
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_67
timestamp 1717613630
transform 0 1 11058 -1 0 22661
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_68
timestamp 1717613630
transform 0 1 10900 -1 0 22573
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_69
timestamp 1717613630
transform 0 1 10742 -1 0 22661
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_70
timestamp 1717613630
transform 0 1 10584 -1 0 22573
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_71
timestamp 1717613630
transform 0 1 10426 -1 0 22225
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_72
timestamp 1717613630
transform 0 1 10268 -1 0 22137
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_73
timestamp 1717613630
transform 0 1 10110 -1 0 22225
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_74
timestamp 1717613630
transform 0 1 9794 -1 0 22225
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_75
timestamp 1717613630
transform 0 1 9952 -1 0 22137
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_76
timestamp 1717613630
transform 0 1 9478 -1 0 22225
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_77
timestamp 1717613630
transform 0 1 9636 -1 0 22137
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_78
timestamp 1717613630
transform 0 1 9162 -1 0 22225
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_79
timestamp 1717613630
transform 0 1 9320 -1 0 22137
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_80
timestamp 1717613630
transform 0 1 8846 -1 0 22661
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_81
timestamp 1717613630
transform 0 1 9004 -1 0 22573
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_82
timestamp 1717613630
transform 0 1 8530 -1 0 22661
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_83
timestamp 1717613630
transform 0 1 8688 -1 0 22573
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_84
timestamp 1717613630
transform 0 1 8688 -1 0 21701
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_85
timestamp 1717613630
transform 0 1 8530 -1 0 21789
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_86
timestamp 1717613630
transform 0 1 9004 -1 0 21701
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_87
timestamp 1717613630
transform 0 1 8846 -1 0 21789
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_88
timestamp 1717613630
transform 0 1 9320 -1 0 21701
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_89
timestamp 1717613630
transform 0 1 9162 -1 0 21789
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_90
timestamp 1717613630
transform 0 1 9636 -1 0 21701
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_91
timestamp 1717613630
transform 0 1 9478 -1 0 21789
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_92
timestamp 1717613630
transform 0 1 9952 -1 0 21701
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_93
timestamp 1717613630
transform 0 1 9794 -1 0 21789
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_94
timestamp 1717613630
transform 0 1 10110 -1 0 21789
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_95
timestamp 1717613630
transform 0 1 10268 -1 0 21701
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_96
timestamp 1717613630
transform 0 1 10426 -1 0 21789
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_97
timestamp 1717613630
transform 0 1 10584 -1 0 21701
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_98
timestamp 1717613630
transform 0 1 10742 -1 0 21789
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_99
timestamp 1717613630
transform 0 1 10900 -1 0 21701
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_100
timestamp 1717613630
transform 0 1 11058 -1 0 21789
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_101
timestamp 1717613630
transform 0 1 11216 -1 0 21701
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_102
timestamp 1717613630
transform 0 1 11374 -1 0 21789
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_103
timestamp 1717613630
transform 0 1 11532 -1 0 21701
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_104
timestamp 1717613630
transform 0 1 11690 -1 0 21789
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_105
timestamp 1717613630
transform 0 1 8846 -1 0 22225
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_106
timestamp 1717613630
transform 0 1 9004 -1 0 22137
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_107
timestamp 1717613630
transform 0 1 8530 -1 0 22225
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_108
timestamp 1717613630
transform 0 1 8688 -1 0 22137
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_109
timestamp 1717613630
transform 0 1 9320 -1 0 22573
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_110
timestamp 1717613630
transform 0 1 9636 -1 0 22573
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_111
timestamp 1717613630
transform 0 1 9952 -1 0 22573
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_112
timestamp 1717613630
transform 0 1 10268 -1 0 22573
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_113
timestamp 1717613630
transform 0 1 9162 -1 0 22661
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_114
timestamp 1717613630
transform 0 1 9478 -1 0 22661
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_115
timestamp 1717613630
transform 0 1 9794 -1 0 22661
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_116
timestamp 1717613630
transform 0 1 10426 -1 0 22661
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_117
timestamp 1717613630
transform 0 1 10110 -1 0 22661
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_118
timestamp 1717613630
transform 0 1 11690 -1 0 22225
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_119
timestamp 1717613630
transform 0 1 11532 -1 0 22137
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_120
timestamp 1717613630
transform 0 1 11374 -1 0 22225
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_121
timestamp 1717613630
transform 0 1 11216 -1 0 22137
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_122
timestamp 1717613630
transform 0 1 11058 -1 0 22225
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_123
timestamp 1717613630
transform 0 1 10900 -1 0 22137
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_124
timestamp 1717613630
transform 0 1 10742 -1 0 22225
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_125
timestamp 1717613630
transform 0 1 10584 -1 0 22137
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_126
timestamp 1717613630
transform 0 1 8688 -1 0 23009
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_127
timestamp 1717613630
transform 0 1 9004 -1 0 23009
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_128
timestamp 1717613630
transform 0 1 9320 -1 0 23009
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_129
timestamp 1717613630
transform 0 1 9636 -1 0 23009
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_130
timestamp 1717613630
transform 0 1 9952 -1 0 23009
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_131
timestamp 1717613630
transform 0 1 10268 -1 0 23009
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_132
timestamp 1717613630
transform 0 1 10584 -1 0 23009
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_133
timestamp 1717613630
transform 0 1 10900 -1 0 23009
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_134
timestamp 1717613630
transform 0 1 11216 -1 0 23009
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_135
timestamp 1717613630
transform 0 1 11532 -1 0 23009
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_136
timestamp 1717613630
transform 0 1 8846 -1 0 23969
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_137
timestamp 1717613630
transform 0 1 8530 -1 0 23969
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_138
timestamp 1717613630
transform 0 1 10426 -1 0 23533
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_139
timestamp 1717613630
transform 0 1 10110 -1 0 23533
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_140
timestamp 1717613630
transform 0 1 9794 -1 0 23533
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_141
timestamp 1717613630
transform 0 1 9478 -1 0 23533
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_142
timestamp 1717613630
transform 0 1 9162 -1 0 23533
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_143
timestamp 1717613630
transform 0 1 11690 -1 0 23969
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_144
timestamp 1717613630
transform 0 1 11374 -1 0 23969
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_145
timestamp 1717613630
transform 0 1 11058 -1 0 23969
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_146
timestamp 1717613630
transform 0 1 10742 -1 0 23969
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_147
timestamp 1717613630
transform 0 1 9004 -1 0 23881
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_148
timestamp 1717613630
transform 0 1 8688 -1 0 23881
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_149
timestamp 1717613630
transform 0 1 8846 -1 0 23097
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_150
timestamp 1717613630
transform 0 1 8530 -1 0 23097
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_151
timestamp 1717613630
transform 0 1 10268 -1 0 23445
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_152
timestamp 1717613630
transform 0 1 9952 -1 0 23445
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_153
timestamp 1717613630
transform 0 1 9636 -1 0 23445
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_154
timestamp 1717613630
transform 0 1 9320 -1 0 23445
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_155
timestamp 1717613630
transform 0 1 10426 -1 0 23097
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_156
timestamp 1717613630
transform 0 1 10110 -1 0 23097
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_157
timestamp 1717613630
transform 0 1 9794 -1 0 23097
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_158
timestamp 1717613630
transform 0 1 9478 -1 0 23097
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_159
timestamp 1717613630
transform 0 1 9162 -1 0 23097
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_160
timestamp 1717613630
transform 0 1 11532 -1 0 23881
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_161
timestamp 1717613630
transform 0 1 11216 -1 0 23881
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_162
timestamp 1717613630
transform 0 1 10900 -1 0 23881
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_163
timestamp 1717613630
transform 0 1 10584 -1 0 23881
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_164
timestamp 1717613630
transform 0 1 11690 -1 0 23097
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_165
timestamp 1717613630
transform 0 1 11374 -1 0 23097
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_166
timestamp 1717613630
transform 0 1 11058 -1 0 23097
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_167
timestamp 1717613630
transform 0 1 10742 -1 0 23097
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_168
timestamp 1717613630
transform 0 1 8846 -1 0 23533
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_169
timestamp 1717613630
transform 0 1 9004 -1 0 23445
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_170
timestamp 1717613630
transform 0 1 8530 -1 0 23533
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_171
timestamp 1717613630
transform 0 1 8688 -1 0 23445
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_172
timestamp 1717613630
transform 0 1 9162 -1 0 23969
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_173
timestamp 1717613630
transform 0 1 9320 -1 0 23881
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_174
timestamp 1717613630
transform 0 1 9794 -1 0 23969
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_175
timestamp 1717613630
transform 0 1 9478 -1 0 23969
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_176
timestamp 1717613630
transform 0 1 9636 -1 0 23881
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_177
timestamp 1717613630
transform 0 1 10110 -1 0 23969
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_178
timestamp 1717613630
transform 0 1 9952 -1 0 23881
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_179
timestamp 1717613630
transform 0 1 10426 -1 0 23969
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_180
timestamp 1717613630
transform 0 1 10268 -1 0 23881
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_181
timestamp 1717613630
transform 0 1 11690 -1 0 23533
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_182
timestamp 1717613630
transform 0 1 11532 -1 0 23445
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_183
timestamp 1717613630
transform 0 1 11374 -1 0 23533
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_184
timestamp 1717613630
transform 0 1 11216 -1 0 23445
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_185
timestamp 1717613630
transform 0 1 11058 -1 0 23533
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_186
timestamp 1717613630
transform 0 1 10900 -1 0 23445
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_187
timestamp 1717613630
transform 0 1 10742 -1 0 23533
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_188
timestamp 1717613630
transform 0 1 10584 -1 0 23445
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_189
timestamp 1717613630
transform 0 1 9004 -1 0 24317
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_190
timestamp 1717613630
transform 0 1 8688 -1 0 24317
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_191
timestamp 1717613630
transform 0 1 8530 -1 0 24405
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_192
timestamp 1717613630
transform 0 1 8846 -1 0 24405
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_193
timestamp 1717613630
transform 0 1 9162 -1 0 24405
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_194
timestamp 1717613630
transform 0 1 9320 -1 0 24317
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_195
timestamp 1717613630
transform 0 1 9794 -1 0 24405
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_196
timestamp 1717613630
transform 0 1 9478 -1 0 24405
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_197
timestamp 1717613630
transform 0 1 9636 -1 0 24317
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_198
timestamp 1717613630
transform 0 1 10110 -1 0 24405
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_199
timestamp 1717613630
transform 0 1 9952 -1 0 24317
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_200
timestamp 1717613630
transform 0 1 10426 -1 0 24405
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_201
timestamp 1717613630
transform 0 1 10268 -1 0 24317
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_202
timestamp 1717613630
transform 0 1 10742 -1 0 24405
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_203
timestamp 1717613630
transform 0 1 10584 -1 0 24317
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_204
timestamp 1717613630
transform 0 1 11058 -1 0 24405
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_205
timestamp 1717613630
transform 0 1 10900 -1 0 24317
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_206
timestamp 1717613630
transform 0 1 11374 -1 0 24405
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_207
timestamp 1717613630
transform 0 1 11216 -1 0 24317
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_208
timestamp 1717613630
transform 0 1 11690 -1 0 24405
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_209
timestamp 1717613630
transform 0 1 11532 -1 0 24317
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_210
timestamp 1717613630
transform 0 1 8846 -1 0 25713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_211
timestamp 1717613630
transform 0 1 9004 -1 0 25625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_212
timestamp 1717613630
transform 0 1 8530 -1 0 25713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_213
timestamp 1717613630
transform 0 1 8688 -1 0 25625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_214
timestamp 1717613630
transform 0 1 10426 -1 0 25277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_215
timestamp 1717613630
transform 0 1 10268 -1 0 25189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_216
timestamp 1717613630
transform 0 1 10110 -1 0 25277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_217
timestamp 1717613630
transform 0 1 9794 -1 0 25277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_218
timestamp 1717613630
transform 0 1 9952 -1 0 25189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_219
timestamp 1717613630
transform 0 1 9478 -1 0 25277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_220
timestamp 1717613630
transform 0 1 9636 -1 0 25189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_221
timestamp 1717613630
transform 0 1 9162 -1 0 25277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_222
timestamp 1717613630
transform 0 1 9320 -1 0 25189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_223
timestamp 1717613630
transform 0 1 11690 -1 0 25713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_224
timestamp 1717613630
transform 0 1 11532 -1 0 25625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_225
timestamp 1717613630
transform 0 1 11374 -1 0 25713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_226
timestamp 1717613630
transform 0 1 11216 -1 0 25625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_227
timestamp 1717613630
transform 0 1 11058 -1 0 25713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_228
timestamp 1717613630
transform 0 1 10900 -1 0 25625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_229
timestamp 1717613630
transform 0 1 10742 -1 0 25713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_230
timestamp 1717613630
transform 0 1 10584 -1 0 25625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_231
timestamp 1717613630
transform 0 1 8846 -1 0 24841
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_232
timestamp 1717613630
transform 0 1 9004 -1 0 24753
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_233
timestamp 1717613630
transform 0 1 8530 -1 0 24841
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_234
timestamp 1717613630
transform 0 1 8688 -1 0 24753
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_235
timestamp 1717613630
transform 0 1 10426 -1 0 24841
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_236
timestamp 1717613630
transform 0 1 10268 -1 0 24753
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_237
timestamp 1717613630
transform 0 1 10110 -1 0 24841
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_238
timestamp 1717613630
transform 0 1 9794 -1 0 24841
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_239
timestamp 1717613630
transform 0 1 9952 -1 0 24753
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_240
timestamp 1717613630
transform 0 1 9478 -1 0 24841
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_241
timestamp 1717613630
transform 0 1 9636 -1 0 24753
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_242
timestamp 1717613630
transform 0 1 9162 -1 0 24841
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_243
timestamp 1717613630
transform 0 1 9320 -1 0 24753
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_244
timestamp 1717613630
transform 0 1 11690 -1 0 24841
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_245
timestamp 1717613630
transform 0 1 11532 -1 0 24753
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_246
timestamp 1717613630
transform 0 1 11374 -1 0 24841
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_247
timestamp 1717613630
transform 0 1 11216 -1 0 24753
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_248
timestamp 1717613630
transform 0 1 11058 -1 0 24841
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_249
timestamp 1717613630
transform 0 1 10900 -1 0 24753
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_250
timestamp 1717613630
transform 0 1 10742 -1 0 24841
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_251
timestamp 1717613630
transform 0 1 10584 -1 0 24753
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_252
timestamp 1717613630
transform 0 1 8846 -1 0 25277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_253
timestamp 1717613630
transform 0 1 9004 -1 0 25189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_254
timestamp 1717613630
transform 0 1 8530 -1 0 25277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_255
timestamp 1717613630
transform 0 1 8688 -1 0 25189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_256
timestamp 1717613630
transform 0 1 9162 -1 0 25713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_257
timestamp 1717613630
transform 0 1 9320 -1 0 25625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_258
timestamp 1717613630
transform 0 1 9478 -1 0 25713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_259
timestamp 1717613630
transform 0 1 9636 -1 0 25625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_260
timestamp 1717613630
transform 0 1 9794 -1 0 25713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_261
timestamp 1717613630
transform 0 1 9952 -1 0 25625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_262
timestamp 1717613630
transform 0 1 10426 -1 0 25713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_263
timestamp 1717613630
transform 0 1 10268 -1 0 25625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_264
timestamp 1717613630
transform 0 1 10110 -1 0 25713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_265
timestamp 1717613630
transform 0 1 11690 -1 0 25277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_266
timestamp 1717613630
transform 0 1 11532 -1 0 25189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_267
timestamp 1717613630
transform 0 1 11374 -1 0 25277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_268
timestamp 1717613630
transform 0 1 11216 -1 0 25189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_269
timestamp 1717613630
transform 0 1 11058 -1 0 25277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_270
timestamp 1717613630
transform 0 1 10900 -1 0 25189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_271
timestamp 1717613630
transform 0 1 10742 -1 0 25277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_272
timestamp 1717613630
transform 0 1 10584 -1 0 25189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_273
timestamp 1717613630
transform 0 1 8846 -1 0 26585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_274
timestamp 1717613630
transform 0 1 9004 -1 0 26497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_275
timestamp 1717613630
transform 0 1 8530 -1 0 26585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_276
timestamp 1717613630
transform 0 1 8688 -1 0 26497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_277
timestamp 1717613630
transform 0 1 10426 -1 0 26585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_278
timestamp 1717613630
transform 0 1 10268 -1 0 26497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_279
timestamp 1717613630
transform 0 1 10110 -1 0 26585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_280
timestamp 1717613630
transform 0 1 9794 -1 0 26585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_281
timestamp 1717613630
transform 0 1 9952 -1 0 26497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_282
timestamp 1717613630
transform 0 1 9478 -1 0 26585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_283
timestamp 1717613630
transform 0 1 9636 -1 0 26497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_284
timestamp 1717613630
transform 0 1 9162 -1 0 26585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_285
timestamp 1717613630
transform 0 1 9320 -1 0 26497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_286
timestamp 1717613630
transform 0 1 11690 -1 0 26585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_287
timestamp 1717613630
transform 0 1 11532 -1 0 26497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_288
timestamp 1717613630
transform 0 1 11374 -1 0 26585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_289
timestamp 1717613630
transform 0 1 11216 -1 0 26497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_290
timestamp 1717613630
transform 0 1 11058 -1 0 26585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_291
timestamp 1717613630
transform 0 1 10900 -1 0 26497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_292
timestamp 1717613630
transform 0 1 10742 -1 0 26585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_293
timestamp 1717613630
transform 0 1 10584 -1 0 26497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_294
timestamp 1717613630
transform 0 1 8846 -1 0 26149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_295
timestamp 1717613630
transform 0 1 9004 -1 0 26061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_296
timestamp 1717613630
transform 0 1 8530 -1 0 26149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_297
timestamp 1717613630
transform 0 1 8688 -1 0 26061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_298
timestamp 1717613630
transform 0 1 10426 -1 0 26149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_299
timestamp 1717613630
transform 0 1 10268 -1 0 26061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_300
timestamp 1717613630
transform 0 1 10110 -1 0 26149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_301
timestamp 1717613630
transform 0 1 9794 -1 0 26149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_302
timestamp 1717613630
transform 0 1 9952 -1 0 26061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_303
timestamp 1717613630
transform 0 1 9478 -1 0 26149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_304
timestamp 1717613630
transform 0 1 9636 -1 0 26061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_305
timestamp 1717613630
transform 0 1 9162 -1 0 26149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_306
timestamp 1717613630
transform 0 1 9320 -1 0 26061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_307
timestamp 1717613630
transform 0 1 11690 -1 0 26149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_308
timestamp 1717613630
transform 0 1 11532 -1 0 26061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_309
timestamp 1717613630
transform 0 1 11374 -1 0 26149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_310
timestamp 1717613630
transform 0 1 11216 -1 0 26061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_311
timestamp 1717613630
transform 0 1 11058 -1 0 26149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_312
timestamp 1717613630
transform 0 1 10900 -1 0 26061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_313
timestamp 1717613630
transform 0 1 10742 -1 0 26149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_314
timestamp 1717613630
transform 0 1 10584 -1 0 26061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_315
timestamp 1717613630
transform 0 1 8688 -1 0 20224
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_316
timestamp 1717613630
transform 0 1 8842 1 0 -12869
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_317
timestamp 1717613630
transform 0 1 8683 1 0 -12777
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_318
timestamp 1717613630
transform 0 1 9737 1 0 -12869
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_319
timestamp 1717613630
transform 0 1 9112 1 0 -13712
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_320
timestamp 1717613630
transform 0 1 9582 1 0 -12777
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_321
timestamp 1717613630
transform 0 1 9266 1 0 -12777
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_322
timestamp 1717613630
transform 0 1 9899 1 0 -12777
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_323
timestamp 1717613630
transform 0 -1 -7377 -1 0 18761
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_324
timestamp 1717613630
transform 0 1 10554 1 0 -13634
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_325
timestamp 1717613630
transform 0 1 8842 1 0 -13638
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_326
timestamp 1717613630
transform 0 1 8683 1 0 -13711
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_327
timestamp 1717613630
transform 0 1 10326 1 0 -12868
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_328
timestamp 1717613630
transform 1 0 -15262 0 -1 -4823
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_329
timestamp 1717613630
transform 0 1 10481 1 0 -12777
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_330
timestamp 1717613630
transform 0 1 10165 1 0 -12777
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_331
timestamp 1717613630
transform 0 1 10798 1 0 -12777
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_332
timestamp 1717613630
transform 0 1 9424 1 0 -12868
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_333
timestamp 1717613630
transform 0 1 11539 1 0 -12869
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_334
timestamp 1717613630
transform 0 1 11226 1 0 -12868
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_335
timestamp 1717613630
transform 0 1 10639 1 0 -12869
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_336
timestamp 1717613630
transform 0 1 11381 1 0 -12777
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_337
timestamp 1717613630
transform 0 1 11065 1 0 -12777
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_338
timestamp 1717613630
transform 0 1 11698 1 0 -12777
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_339
timestamp 1717613630
transform 0 1 9272 1 0 -13636
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_340
timestamp 1717613630
transform 0 1 10133 1 0 -14503
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_341
timestamp 1717613630
transform 0 1 9862 1 0 -13636
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_342
timestamp 1717613630
transform 0 1 11037 1 0 -13637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_343
timestamp 1717613630
transform 0 1 10289 1 0 -13710
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_344
timestamp 1717613630
transform 0 1 10799 1 0 -13711
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_345
timestamp 1717613630
transform 0 1 9541 1 0 -13636
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_346
timestamp 1717613630
transform 0 1 9861 1 0 -14433
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_347
timestamp 1717613630
transform 0 1 9545 1 0 -14433
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_348
timestamp 1717613630
transform 0 1 9229 1 0 -14433
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_349
timestamp 1717613630
transform 0 1 9388 1 0 -14507
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_350
timestamp 1717613630
transform 1 0 -15591 0 -1 -6473
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_351
timestamp 1717613630
transform 0 1 10860 1 0 -14584
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_352
timestamp 1717613630
transform 1 0 -13970 0 -1 -4935
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_353
timestamp 1717613630
transform 1 0 -13967 0 -1 -5086
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_354
timestamp 1717613630
transform 0 1 9702 1 0 -13711
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_355
timestamp 1717613630
transform 0 1 11307 1 0 -13638
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_356
timestamp 1717613630
transform 0 1 10132 1 0 -13710
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_357
timestamp 1717613630
transform 0 1 11623 1 0 -13638
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_358
timestamp 1717613630
transform 0 1 11468 1 0 -13707
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_359
timestamp 1717613630
transform 1 0 -13383 0 -1 -6391
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_360
timestamp 1717613630
transform 1 0 -13856 0 -1 -6632
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_361
timestamp 1717613630
transform 0 1 10993 1 0 -14434
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_362
timestamp 1717613630
transform 0 1 11152 1 0 -14508
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_363
timestamp 1717613630
transform 0 1 11309 1 0 -14434
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_364
timestamp 1717613630
transform 0 1 11467 1 0 -14508
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_365
timestamp 1717613630
transform 0 1 11625 1 0 -14434
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_366
timestamp 1717613630
transform 0 1 9703 1 0 -14507
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_367
timestamp 1717613630
transform 1 0 -15376 0 -1 -6632
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_368
timestamp 1717613630
transform 0 -1 -7295 -1 0 18941
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_369
timestamp 1717613630
transform 0 1 10564 1 0 -14433
box 16088 -7932 16222 -7868
use sky130_fd_pr__nfet_g5v0d10v5_FJGQFC  XM1 paramcells
timestamp 1717692607
transform 1 0 1801 0 1 2481
box -357 -358 357 358
use sky130_fd_pr__pfet_g5v0d10v5_KLWMS5  XM5 paramcells
timestamp 1717691772
transform 1 0 2583 0 1 3332
box -545 -397 545 397
use sky130_fd_pr__pfet_g5v0d10v5_KLWMS5  XM6
timestamp 1717691772
transform 1 0 3483 0 1 3332
box -545 -397 545 397
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM7 paramcells
timestamp 1717690002
transform 1 0 3567 0 1 2481
box -357 -358 357 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQFS  XM8 paramcells
timestamp 1717691772
transform 1 0 2310 0 1 2481
box -278 -358 278 358
use sky130_fd_pr__nfet_05v0_nvt_BH6ZTK  XM9 paramcells
timestamp 1717692607
transform 1 0 2899 0 1 2481
box -437 -358 437 358
use sky130_fd_pr__nfet_g5v0d10v5_H7BQFY  XM10 paramcells
timestamp 1717691772
transform 1 0 1645 0 1 1685
box -515 -358 515 358
use sky130_fd_pr__pfet_g5v0d10v5_AQ2WAW  XM12 paramcells
timestamp 1717690002
transform 1 0 2210 0 1 4113
box -1809 -397 1809 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQFS  XM13
timestamp 1717691772
transform 1 0 2312 0 1 1685
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_Z8JNCQ  XM20 paramcells
timestamp 1717691772
transform 1 0 2210 0 1 7551
box -1809 -3231 1809 3231
use sky130_fd_pr__nfet_g5v0d10v5_H7BQ24  XM22 paramcells
timestamp 1717690002
transform 1 0 3409 0 1 1684
box -515 -358 515 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQFS  XM24
timestamp 1717691772
transform 1 0 2742 0 1 1685
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_KLJMY6  XM25 paramcells
timestamp 1717692607
transform 1 0 862 0 1 3332
box -466 -397 466 397
use sky130_fd_pr__pfet_g5v0d10v5_KLWMS5  XM27
timestamp 1717691772
transform 1 0 1683 0 1 3332
box -545 -397 545 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQFS  XM29
timestamp 1717691772
transform 1 0 1292 0 1 2481
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQFS  XM30
timestamp 1717691772
transform 1 0 862 0 1 2481
box -278 -358 278 358
use sky130_fd_pr__res_xhigh_po_0p35_HLA228  XR1 paramcells
timestamp 1717716768
transform 0 1 2187 -1 0 807
box -367 -1748 367 1748
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XXD1 paramcells
timestamp 1717690002
transform 1 0 771 0 1 1552
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XXD2
timestamp 1717690002
transform 1 0 771 0 1 1812
box -183 -183 183 183
<< labels >>
flabel metal2 276 10482 476 10682 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal2 3906 4358 4106 4558 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal2 1171 3244 1171 3244 0 FreeSans 400 0 0 0 vcomp
flabel metal2 257 2980 457 3180 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal2 2021 1563 2021 1563 0 FreeSans 400 0 0 0 nbias
flabel metal2 283 1975 483 2175 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal2 261 1247 461 1447 0 FreeSans 256 0 0 0 ena
port 2 nsew
flabel metal1 704 2881 704 2881 0 FreeSans 400 90 0 0 pbias
flabel metal1 0 0 108 149 0 FreeSans 960 0 0 0 vsub
port 5 nsew
<< end >>
