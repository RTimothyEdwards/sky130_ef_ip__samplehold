magic
tech sky130A
magscale 1 2
timestamp 1717718523
<< dnwell >>
rect 3092 -5410 7008 5247
<< nwell >>
rect 2983 5041 7117 5356
rect 2983 -5204 3298 5041
rect 6802 -5204 7117 5041
rect 2983 -5519 7117 -5204
<< mvpsubdiff >>
rect 2863 5453 2923 5487
rect 7179 5453 7239 5487
rect 2863 5427 2897 5453
rect 7205 5427 7239 5453
rect 2863 -5606 2897 -5510
rect 7205 -5606 7239 -5510
rect 2863 -5640 2923 -5606
rect 7179 -5640 7239 -5606
<< mvnsubdiff >>
rect 3049 5270 7051 5290
rect 3049 5236 3129 5270
rect 6971 5236 7051 5270
rect 3049 5216 7051 5236
rect 3049 5210 3123 5216
rect 3049 -5373 3069 5210
rect 3103 -5373 3123 5210
rect 3049 -5379 3123 -5373
rect 6977 5210 7051 5216
rect 6977 -5373 6997 5210
rect 7031 -5373 7051 5210
rect 6977 -5379 7051 -5373
rect 3049 -5399 7051 -5379
rect 3049 -5433 3129 -5399
rect 6971 -5433 7051 -5399
rect 3049 -5453 7051 -5433
<< mvpsubdiffcont >>
rect 2923 5453 7179 5487
rect 2863 -5510 2897 5427
rect 7205 -5510 7239 5427
rect 2923 -5640 7179 -5606
<< mvnsubdiffcont >>
rect 3129 5236 6971 5270
rect 3069 -5373 3103 5210
rect 6997 -5373 7031 5210
rect 3129 -5433 6971 -5399
<< locali >>
rect 2863 5487 7240 5489
rect 2863 5453 2923 5487
rect 7179 5453 7240 5487
rect 2863 5431 3027 5453
rect 2863 5427 2908 5431
rect 2897 -5429 2908 5427
rect 2952 5409 3027 5431
rect 7091 5438 7240 5453
rect 7091 5409 7164 5438
rect 7210 5427 7240 5438
rect 2952 5389 7164 5409
rect 2952 -5429 2971 5389
rect 2897 -5510 2971 -5429
rect 3042 5299 3146 5303
rect 3042 5280 7051 5299
rect 3042 5270 3144 5280
rect 6946 5270 7051 5280
rect 3042 5236 3129 5270
rect 6971 5236 7051 5270
rect 3042 5228 3144 5236
rect 6946 5228 7051 5236
rect 3042 5210 7051 5228
rect 3042 5200 3069 5210
rect 3103 5208 6997 5210
rect 3103 5200 3146 5208
rect 3042 -5348 3065 5200
rect 3110 -5348 3146 5200
rect 6950 5187 6997 5208
rect 3235 5066 6836 5092
rect 3235 5031 3384 5066
rect 6633 5063 6836 5066
rect 6633 5031 6793 5063
rect 3235 5003 6793 5031
rect 3235 4770 3405 5003
rect 3235 -1823 3246 4770
rect 3300 -1168 3405 4770
rect 6747 -1168 6793 5003
rect 3300 -1200 6793 -1168
rect 3300 -1242 3509 -1200
rect 6653 -1242 6793 -1200
rect 3300 -1269 6793 -1242
rect 3300 -1783 3405 -1269
rect 6747 -1783 6793 -1269
rect 3300 -1799 6793 -1783
rect 3300 -1823 3540 -1799
rect 3235 -1834 3540 -1823
rect 5787 -1801 6793 -1799
rect 5787 -1834 5977 -1801
rect 3235 -1835 5977 -1834
rect 6669 -1835 6793 -1801
rect 3235 -1872 6793 -1835
rect 3290 -1974 6793 -1944
rect 3290 -1975 5095 -1974
rect 3290 -2023 3338 -1975
rect 4871 -2021 5095 -1975
rect 5809 -1978 6793 -1974
rect 5809 -2021 5986 -1978
rect 4871 -2023 5986 -2021
rect 3290 -2025 5986 -2023
rect 6662 -2025 6793 -1978
rect 3290 -2055 6793 -2025
rect 3311 -2550 3422 -2055
rect 6743 -2512 6793 -2055
rect 6832 -1872 6836 5063
rect 6832 -1945 6842 -1944
rect 6832 -2512 6854 -1945
rect 6743 -2550 6854 -2512
rect 3302 -2661 6854 -2550
rect 6950 -2558 6987 5187
rect 6950 -2585 6997 -2558
rect 3458 -2836 6768 -2813
rect 3458 -2921 6687 -2836
rect 3458 -3389 3566 -2921
rect 6660 -3389 6687 -2921
rect 3457 -3419 6687 -3389
rect 3457 -3470 3727 -3419
rect 5077 -3444 6687 -3419
rect 6742 -3444 6768 -2836
rect 5077 -3470 6768 -3444
rect 3457 -3497 6768 -3470
rect 4056 -3612 6768 -3608
rect 3449 -3640 6768 -3612
rect 3449 -3677 3597 -3640
rect 5605 -3653 6768 -3640
rect 5605 -3677 6688 -3653
rect 3449 -3693 6688 -3677
rect 3449 -4192 3550 -3693
rect 3756 -3717 6688 -3693
rect 3756 -4132 3798 -3717
rect 3755 -4192 3798 -4132
rect 3449 -4197 3798 -4192
rect 3836 -3722 6688 -3717
rect 3836 -3730 4056 -3722
rect 3836 -4197 3973 -3730
rect 3449 -4198 3973 -4197
rect 4014 -4192 4056 -3730
rect 5389 -4192 5517 -3854
rect 6654 -4192 6688 -3722
rect 4014 -4198 6688 -4192
rect 3449 -4221 6688 -4198
rect 3449 -4269 4160 -4221
rect 5053 -4261 6688 -4221
rect 6743 -4261 6768 -3653
rect 5053 -4269 6768 -4261
rect 3449 -4306 6768 -4269
rect 3755 -4437 4056 -4306
rect 3305 -4457 6878 -4437
rect 3305 -4471 6823 -4457
rect 3305 -4507 3427 -4471
rect 6153 -4507 6823 -4471
rect 3305 -4545 6823 -4507
rect 3305 -4898 3400 -4545
rect 3305 -5043 3322 -4898
rect 3369 -5043 3400 -4898
rect 3305 -5092 3400 -5043
rect 6744 -5092 6823 -4545
rect 3305 -5121 6823 -5092
rect 6863 -5121 6878 -4457
rect 3305 -5124 6878 -5121
rect 3305 -5161 3317 -5124
rect 6782 -5161 6878 -5124
rect 3305 -5198 6878 -5161
rect 3042 -5373 3069 -5348
rect 3103 -5359 3146 -5348
rect 3103 -5373 6997 -5359
rect 7031 -2585 7051 5210
rect 7031 -5373 7058 -5359
rect 3042 -5387 7058 -5373
rect 3042 -5441 3118 -5387
rect 6980 -5441 7058 -5387
rect 3042 -5471 7058 -5441
rect 2863 -5538 2971 -5510
rect 7141 -5538 7164 5389
rect 7239 -5510 7240 5427
rect 2863 -5568 7164 -5538
rect 2863 -5606 3011 -5568
rect 7122 -5570 7164 -5568
rect 7210 -5570 7240 -5510
rect 7122 -5606 7240 -5570
rect 2863 -5640 2923 -5606
rect 7179 -5640 7240 -5606
<< viali >>
rect 3027 5453 7091 5455
rect 2908 -5429 2952 5431
rect 3027 5409 7091 5453
rect 7164 5427 7210 5438
rect 3144 5270 6946 5280
rect 3144 5236 6946 5270
rect 3144 5228 6946 5236
rect 3065 -5348 3069 5200
rect 3069 -5348 3103 5200
rect 3103 -5348 3110 5200
rect 3384 5031 6633 5066
rect 3246 -1823 3300 4770
rect 3509 -1242 6653 -1200
rect 3540 -1834 5787 -1799
rect 5977 -1835 6669 -1801
rect 3338 -2023 4871 -1975
rect 5095 -2021 5809 -1974
rect 5986 -2025 6662 -1978
rect 6793 -2512 6832 5063
rect 6987 -2558 6997 5187
rect 6997 -2558 7030 5187
rect 3727 -3470 5077 -3419
rect 6687 -3444 6742 -2836
rect 3597 -3677 5605 -3640
rect 3798 -4197 3836 -3717
rect 3973 -4198 4014 -3730
rect 4160 -4269 5053 -4221
rect 6688 -4261 6743 -3653
rect 3427 -4507 6153 -4471
rect 3322 -5043 3369 -4898
rect 6823 -5121 6863 -4457
rect 3317 -5161 6782 -5124
rect 3118 -5399 6980 -5387
rect 3118 -5433 3129 -5399
rect 3129 -5433 6971 -5399
rect 6971 -5433 6980 -5399
rect 3118 -5441 6980 -5433
rect 7164 -5510 7205 5427
rect 7205 -5510 7210 5427
rect 3011 -5606 7122 -5568
rect 7164 -5570 7210 -5510
rect 3011 -5614 7122 -5606
<< metal1 >>
rect 2863 5455 7240 5489
rect 2863 5431 3027 5455
rect 2863 -5429 2908 5431
rect 2952 5409 3027 5431
rect 7091 5438 7240 5455
rect 7091 5409 7164 5438
rect 2952 5389 7164 5409
rect 2952 -5429 2971 5389
rect 2863 -5538 2971 -5429
rect 3042 5299 3146 5303
rect 3042 5280 7051 5299
rect 3042 5228 3144 5280
rect 6946 5228 7051 5280
rect 3042 5208 7051 5228
rect 3042 5200 3146 5208
rect 3042 -5348 3065 5200
rect 3110 -1147 3146 5200
rect 3216 5093 3321 5208
rect 6770 5094 6875 5208
rect 6950 5187 7051 5208
rect 6770 5093 6877 5094
rect 3216 5092 6877 5093
rect 3213 5078 6877 5092
rect 3213 5066 3407 5078
rect 6621 5066 6877 5078
rect 3213 5031 3384 5066
rect 6633 5063 6877 5066
rect 6633 5031 6793 5063
rect 3213 5024 3407 5031
rect 6621 5024 6793 5031
rect 3213 5004 6793 5024
rect 3213 4788 3320 5004
rect 3213 -1147 3223 4788
rect 3110 -1265 3223 -1147
rect 3110 -1947 3146 -1265
rect 3213 -1947 3223 -1265
rect 3110 -2056 3223 -1947
rect 3110 -5348 3146 -2056
rect 3213 -2255 3223 -2056
rect 3309 -1969 3320 4788
rect 3368 4928 3534 4932
rect 3713 4928 3745 4932
rect 3871 4928 3903 4932
rect 4029 4928 4061 4932
rect 4187 4928 4219 4932
rect 4345 4928 4377 4932
rect 4503 4928 4535 4932
rect 4661 4928 4693 4932
rect 4819 4928 4851 4932
rect 4977 4928 5009 4932
rect 5135 4928 5167 4932
rect 5293 4928 5325 4932
rect 5451 4928 5483 4932
rect 5609 4928 5641 4932
rect 5767 4928 5799 4932
rect 5925 4928 5957 4932
rect 6083 4928 6115 4932
rect 6241 4928 6273 4932
rect 6399 4928 6431 4932
rect 6557 4928 6589 4932
rect 3368 4891 6628 4928
rect 3368 4886 3534 4891
rect 3368 4604 3415 4886
rect 3368 4600 3534 4604
rect 3555 4600 3587 4891
rect 3713 4600 3745 4891
rect 3871 4600 3903 4891
rect 4029 4600 4061 4891
rect 4187 4600 4219 4891
rect 4345 4600 4377 4891
rect 4503 4600 4535 4891
rect 4661 4600 4693 4891
rect 4819 4600 4851 4891
rect 4977 4600 5009 4891
rect 5135 4600 5167 4891
rect 5293 4600 5325 4891
rect 5451 4600 5483 4891
rect 5609 4600 5641 4891
rect 5767 4600 5799 4891
rect 5925 4600 5957 4891
rect 6083 4600 6115 4891
rect 6241 4600 6273 4891
rect 6399 4600 6431 4891
rect 6557 4600 6589 4891
rect 3368 4563 6620 4600
rect 3368 4558 3534 4563
rect 3368 4496 3415 4558
rect 3368 4492 3534 4496
rect 3555 4492 3587 4563
rect 3713 4492 3745 4563
rect 3871 4492 3903 4563
rect 4029 4492 4061 4563
rect 4187 4492 4219 4563
rect 4345 4492 4377 4563
rect 4503 4492 4535 4563
rect 4661 4492 4693 4563
rect 4819 4492 4851 4563
rect 4977 4492 5009 4563
rect 5135 4492 5167 4563
rect 5293 4492 5325 4563
rect 5451 4492 5483 4563
rect 5609 4492 5641 4563
rect 5767 4492 5799 4563
rect 5925 4492 5957 4563
rect 6083 4492 6115 4563
rect 6241 4492 6273 4563
rect 6399 4492 6431 4563
rect 6557 4492 6589 4563
rect 3368 4455 6628 4492
rect 3368 4450 3534 4455
rect 3368 4168 3415 4450
rect 3368 4164 3534 4168
rect 3555 4164 3587 4455
rect 3713 4164 3745 4455
rect 3871 4164 3903 4455
rect 4029 4164 4061 4455
rect 4187 4164 4219 4455
rect 4345 4164 4377 4455
rect 4503 4164 4535 4455
rect 4661 4164 4693 4455
rect 4819 4164 4851 4455
rect 4977 4164 5009 4455
rect 5135 4164 5167 4455
rect 5293 4164 5325 4455
rect 5451 4164 5483 4455
rect 5609 4164 5641 4455
rect 5767 4164 5799 4455
rect 5925 4164 5957 4455
rect 6083 4164 6115 4455
rect 6241 4164 6273 4455
rect 6399 4164 6431 4455
rect 6557 4164 6589 4455
rect 3368 4127 6620 4164
rect 3368 4122 3534 4127
rect 3368 4060 3415 4122
rect 3368 4056 3534 4060
rect 3555 4056 3587 4127
rect 3713 4056 3745 4127
rect 3871 4056 3903 4127
rect 4029 4056 4061 4127
rect 4187 4056 4219 4127
rect 4345 4056 4377 4127
rect 4503 4056 4535 4127
rect 4661 4056 4693 4127
rect 4819 4056 4851 4127
rect 4977 4056 5009 4127
rect 5135 4056 5167 4127
rect 5293 4056 5325 4127
rect 5451 4056 5483 4127
rect 5609 4056 5641 4127
rect 5767 4056 5799 4127
rect 5925 4056 5957 4127
rect 6083 4056 6115 4127
rect 6241 4056 6273 4127
rect 6399 4056 6431 4127
rect 6557 4056 6589 4127
rect 3368 4019 6628 4056
rect 3368 4014 3534 4019
rect 3368 3732 3415 4014
rect 3368 3728 3534 3732
rect 3555 3728 3587 4019
rect 3713 3728 3745 4019
rect 3871 3728 3903 4019
rect 4029 3728 4061 4019
rect 4187 3728 4219 4019
rect 4345 3728 4377 4019
rect 4503 3728 4535 4019
rect 4661 3728 4693 4019
rect 4819 3728 4851 4019
rect 4977 3728 5009 4019
rect 5135 3728 5167 4019
rect 5293 3728 5325 4019
rect 5451 3728 5483 4019
rect 5609 3728 5641 4019
rect 5767 3728 5799 4019
rect 5925 3728 5957 4019
rect 6083 3728 6115 4019
rect 6241 3728 6273 4019
rect 6399 3728 6431 4019
rect 6557 3728 6589 4019
rect 3368 3691 6620 3728
rect 3368 3686 3534 3691
rect 3368 3624 3415 3686
rect 3368 3620 3534 3624
rect 3555 3620 3587 3691
rect 3713 3620 3745 3691
rect 3871 3620 3903 3691
rect 4029 3620 4061 3691
rect 4187 3620 4219 3691
rect 4345 3620 4377 3691
rect 4503 3620 4535 3691
rect 4661 3620 4693 3691
rect 4819 3620 4851 3691
rect 4977 3620 5009 3691
rect 5135 3620 5167 3691
rect 5293 3620 5325 3691
rect 5451 3620 5483 3691
rect 5609 3620 5641 3691
rect 5767 3620 5799 3691
rect 5925 3620 5957 3691
rect 6083 3620 6115 3691
rect 6241 3620 6273 3691
rect 6399 3620 6431 3691
rect 6557 3620 6589 3691
rect 3368 3583 6628 3620
rect 3368 3578 3534 3583
rect 3368 3296 3415 3578
rect 3368 3292 3534 3296
rect 3555 3292 3587 3583
rect 3713 3292 3745 3583
rect 3871 3292 3903 3583
rect 4029 3292 4061 3583
rect 4187 3292 4219 3583
rect 4345 3292 4377 3583
rect 4503 3292 4535 3583
rect 4661 3292 4693 3583
rect 4819 3292 4851 3583
rect 4977 3292 5009 3583
rect 5135 3292 5167 3583
rect 5293 3292 5325 3583
rect 5451 3292 5483 3583
rect 5609 3292 5641 3583
rect 5767 3292 5799 3583
rect 5925 3292 5957 3583
rect 6083 3292 6115 3583
rect 6241 3292 6273 3583
rect 6399 3292 6431 3583
rect 6557 3292 6589 3583
rect 3368 3255 6620 3292
rect 3368 3250 3534 3255
rect 3368 3188 3415 3250
rect 3368 3184 3534 3188
rect 3555 3184 3587 3255
rect 3713 3184 3745 3255
rect 3871 3184 3903 3255
rect 4029 3184 4061 3255
rect 4187 3184 4219 3255
rect 4345 3184 4377 3255
rect 4503 3184 4535 3255
rect 4661 3184 4693 3255
rect 4819 3184 4851 3255
rect 4977 3184 5009 3255
rect 5135 3184 5167 3255
rect 5293 3184 5325 3255
rect 5451 3184 5483 3255
rect 5609 3184 5641 3255
rect 5767 3184 5799 3255
rect 5925 3184 5957 3255
rect 6083 3184 6115 3255
rect 6241 3184 6273 3255
rect 6399 3184 6431 3255
rect 6557 3184 6589 3255
rect 3368 3147 6628 3184
rect 3368 3142 3534 3147
rect 3368 2860 3415 3142
rect 3368 2856 3534 2860
rect 3555 2856 3587 3147
rect 3713 2856 3745 3147
rect 3871 2856 3903 3147
rect 4029 2856 4061 3147
rect 4187 2856 4219 3147
rect 4345 2856 4377 3147
rect 4503 2856 4535 3147
rect 4661 2856 4693 3147
rect 4819 2856 4851 3147
rect 4977 2856 5009 3147
rect 5135 2856 5167 3147
rect 5293 2856 5325 3147
rect 5451 2856 5483 3147
rect 5609 2856 5641 3147
rect 5767 2856 5799 3147
rect 5925 2856 5957 3147
rect 6083 2856 6115 3147
rect 6241 2856 6273 3147
rect 6399 2856 6431 3147
rect 6557 2856 6589 3147
rect 3368 2819 6620 2856
rect 3368 2814 3534 2819
rect 3368 2752 3415 2814
rect 3368 2748 3534 2752
rect 3555 2748 3587 2819
rect 3713 2748 3745 2819
rect 3871 2748 3903 2819
rect 4029 2748 4061 2819
rect 4187 2748 4219 2819
rect 4345 2748 4377 2819
rect 4503 2748 4535 2819
rect 4661 2748 4693 2819
rect 4819 2748 4851 2819
rect 4977 2748 5009 2819
rect 5135 2748 5167 2819
rect 5293 2748 5325 2819
rect 5451 2748 5483 2819
rect 5609 2748 5641 2819
rect 5767 2748 5799 2819
rect 5925 2748 5957 2819
rect 6083 2748 6115 2819
rect 6241 2748 6273 2819
rect 6399 2748 6431 2819
rect 6557 2748 6589 2819
rect 3368 2711 6628 2748
rect 3368 2706 3534 2711
rect 3368 2424 3415 2706
rect 3368 2420 3534 2424
rect 3555 2420 3587 2711
rect 3713 2420 3745 2711
rect 3871 2420 3903 2711
rect 4029 2420 4061 2711
rect 4187 2420 4219 2711
rect 4345 2420 4377 2711
rect 4503 2420 4535 2711
rect 4661 2420 4693 2711
rect 4819 2420 4851 2711
rect 4977 2420 5009 2711
rect 5135 2420 5167 2711
rect 5293 2420 5325 2711
rect 5451 2420 5483 2711
rect 5609 2420 5641 2711
rect 5767 2420 5799 2711
rect 5925 2420 5957 2711
rect 6083 2420 6115 2711
rect 6241 2420 6273 2711
rect 6399 2420 6431 2711
rect 6557 2420 6589 2711
rect 3368 2383 6620 2420
rect 3368 2378 3534 2383
rect 3368 2316 3415 2378
rect 3368 2312 3534 2316
rect 3555 2312 3587 2383
rect 3713 2312 3745 2383
rect 3871 2312 3903 2383
rect 4029 2312 4061 2383
rect 4187 2312 4219 2383
rect 4345 2312 4377 2383
rect 4503 2312 4535 2383
rect 4661 2312 4693 2383
rect 4819 2312 4851 2383
rect 4977 2312 5009 2383
rect 5135 2312 5167 2383
rect 5293 2312 5325 2383
rect 5451 2312 5483 2383
rect 5609 2312 5641 2383
rect 5767 2312 5799 2383
rect 5925 2312 5957 2383
rect 6083 2312 6115 2383
rect 6241 2312 6273 2383
rect 6399 2312 6431 2383
rect 6557 2312 6589 2383
rect 3368 2275 6628 2312
rect 3368 2270 3534 2275
rect 3368 1988 3415 2270
rect 3368 1984 3534 1988
rect 3555 1984 3587 2275
rect 3713 1984 3745 2275
rect 3871 1984 3903 2275
rect 4029 1984 4061 2275
rect 4187 1984 4219 2275
rect 4345 1984 4377 2275
rect 4503 1984 4535 2275
rect 4661 1984 4693 2275
rect 4819 1984 4851 2275
rect 4977 1984 5009 2275
rect 5135 1984 5167 2275
rect 5293 1984 5325 2275
rect 5451 1984 5483 2275
rect 5609 1984 5641 2275
rect 5767 1984 5799 2275
rect 5925 1984 5957 2275
rect 6083 1984 6115 2275
rect 6241 1984 6273 2275
rect 6399 1984 6431 2275
rect 6557 1984 6589 2275
rect 3368 1947 6620 1984
rect 3368 1942 3534 1947
rect 3368 1880 3415 1942
rect 3368 1876 3534 1880
rect 3555 1876 3587 1947
rect 3713 1876 3745 1947
rect 3871 1876 3903 1947
rect 4029 1876 4061 1947
rect 4187 1876 4219 1947
rect 4345 1876 4377 1947
rect 4503 1876 4535 1947
rect 4661 1876 4693 1947
rect 4819 1876 4851 1947
rect 4977 1876 5009 1947
rect 5135 1876 5167 1947
rect 5293 1876 5325 1947
rect 5451 1876 5483 1947
rect 5609 1876 5641 1947
rect 5767 1876 5799 1947
rect 5925 1876 5957 1947
rect 6083 1876 6115 1947
rect 6241 1876 6273 1947
rect 6399 1876 6431 1947
rect 6557 1876 6589 1947
rect 3368 1839 6628 1876
rect 3368 1834 3534 1839
rect 3368 1552 3415 1834
rect 3368 1548 3534 1552
rect 3555 1548 3587 1839
rect 3713 1548 3745 1839
rect 3871 1548 3903 1839
rect 4029 1548 4061 1839
rect 4187 1548 4219 1839
rect 4345 1548 4377 1839
rect 4503 1548 4535 1839
rect 4661 1548 4693 1839
rect 4819 1548 4851 1839
rect 4977 1548 5009 1839
rect 5135 1548 5167 1839
rect 5293 1548 5325 1839
rect 5451 1548 5483 1839
rect 5609 1548 5641 1839
rect 5767 1548 5799 1839
rect 5925 1548 5957 1839
rect 6083 1548 6115 1839
rect 6241 1548 6273 1839
rect 6399 1548 6431 1839
rect 6557 1548 6589 1839
rect 3368 1511 6620 1548
rect 3368 1506 3534 1511
rect 3368 1444 3415 1506
rect 3368 1440 3534 1444
rect 3555 1440 3587 1511
rect 3713 1440 3745 1511
rect 3871 1440 3903 1511
rect 4029 1440 4061 1511
rect 4187 1440 4219 1511
rect 4345 1440 4377 1511
rect 4503 1440 4535 1511
rect 4661 1440 4693 1511
rect 4819 1440 4851 1511
rect 4977 1440 5009 1511
rect 5135 1440 5167 1511
rect 5293 1440 5325 1511
rect 5451 1440 5483 1511
rect 5609 1440 5641 1511
rect 5767 1440 5799 1511
rect 5925 1440 5957 1511
rect 6083 1440 6115 1511
rect 6241 1440 6273 1511
rect 6399 1440 6431 1511
rect 6557 1440 6589 1511
rect 3368 1403 6628 1440
rect 3368 1398 3534 1403
rect 3368 1116 3415 1398
rect 3368 1112 3534 1116
rect 3555 1112 3587 1403
rect 3713 1112 3745 1403
rect 3871 1112 3903 1403
rect 4029 1112 4061 1403
rect 4187 1112 4219 1403
rect 4345 1112 4377 1403
rect 4503 1112 4535 1403
rect 4661 1112 4693 1403
rect 4819 1112 4851 1403
rect 4977 1112 5009 1403
rect 5135 1112 5167 1403
rect 5293 1112 5325 1403
rect 5451 1112 5483 1403
rect 5609 1112 5641 1403
rect 5767 1112 5799 1403
rect 5925 1112 5957 1403
rect 6083 1112 6115 1403
rect 6241 1112 6273 1403
rect 6399 1112 6431 1403
rect 6557 1112 6589 1403
rect 3368 1075 6620 1112
rect 3368 1070 3534 1075
rect 3368 1008 3415 1070
rect 3368 1004 3534 1008
rect 3555 1004 3587 1075
rect 3713 1004 3745 1075
rect 3871 1004 3903 1075
rect 4029 1004 4061 1075
rect 4187 1004 4219 1075
rect 4345 1004 4377 1075
rect 4503 1004 4535 1075
rect 4661 1004 4693 1075
rect 4819 1004 4851 1075
rect 4977 1004 5009 1075
rect 5135 1004 5167 1075
rect 5293 1004 5325 1075
rect 5451 1004 5483 1075
rect 5609 1004 5641 1075
rect 5767 1004 5799 1075
rect 5925 1004 5957 1075
rect 6083 1004 6115 1075
rect 6241 1004 6273 1075
rect 6399 1004 6431 1075
rect 6557 1004 6589 1075
rect 3368 967 6628 1004
rect 3368 962 3534 967
rect 3368 680 3415 962
rect 3368 676 3534 680
rect 3555 676 3587 967
rect 3713 676 3745 967
rect 3871 676 3903 967
rect 4029 676 4061 967
rect 4187 676 4219 967
rect 4345 676 4377 967
rect 4503 676 4535 967
rect 4661 676 4693 967
rect 4819 676 4851 967
rect 4977 676 5009 967
rect 5135 676 5167 967
rect 5293 676 5325 967
rect 5451 676 5483 967
rect 5609 676 5641 967
rect 5767 676 5799 967
rect 5925 676 5957 967
rect 6083 676 6115 967
rect 6241 676 6273 967
rect 6399 676 6431 967
rect 6557 676 6589 967
rect 3368 639 6620 676
rect 3368 634 3534 639
rect 3368 572 3415 634
rect 3368 568 3534 572
rect 3555 568 3587 639
rect 3713 568 3745 639
rect 3871 568 3903 639
rect 4029 568 4061 639
rect 4187 568 4219 639
rect 4345 568 4377 639
rect 4503 568 4535 639
rect 4661 568 4693 639
rect 4819 568 4851 639
rect 4977 568 5009 639
rect 5135 568 5167 639
rect 5293 568 5325 639
rect 5451 568 5483 639
rect 5609 568 5641 639
rect 5767 568 5799 639
rect 5925 568 5957 639
rect 6083 568 6115 639
rect 6241 568 6273 639
rect 6399 568 6431 639
rect 6557 568 6589 639
rect 3368 531 6628 568
rect 3368 526 3534 531
rect 3368 244 3415 526
rect 3368 240 3534 244
rect 3555 240 3587 531
rect 3713 240 3745 531
rect 3871 240 3903 531
rect 4029 240 4061 531
rect 4187 240 4219 531
rect 4345 240 4377 531
rect 4503 240 4535 531
rect 4661 240 4693 531
rect 4819 240 4851 531
rect 4977 240 5009 531
rect 5135 240 5167 531
rect 5293 240 5325 531
rect 5451 240 5483 531
rect 5609 240 5641 531
rect 5767 240 5799 531
rect 5925 240 5957 531
rect 6083 240 6115 531
rect 6241 240 6273 531
rect 6399 240 6431 531
rect 6557 240 6589 531
rect 3368 203 6620 240
rect 3368 198 3534 203
rect 3368 136 3415 198
rect 3368 132 3534 136
rect 3555 132 3587 203
rect 3713 132 3745 203
rect 3871 132 3903 203
rect 4029 132 4061 203
rect 4187 132 4219 203
rect 4345 132 4377 203
rect 4503 132 4535 203
rect 4661 132 4693 203
rect 4819 132 4851 203
rect 4977 132 5009 203
rect 5135 132 5167 203
rect 5293 132 5325 203
rect 5451 132 5483 203
rect 5609 132 5641 203
rect 5767 132 5799 203
rect 5925 132 5957 203
rect 6083 132 6115 203
rect 6241 132 6273 203
rect 6399 132 6431 203
rect 6557 132 6589 203
rect 3368 95 6628 132
rect 3368 90 3534 95
rect 3368 -192 3415 90
rect 3368 -196 3534 -192
rect 3555 -196 3587 95
rect 3713 -196 3745 95
rect 3871 -196 3903 95
rect 4029 -196 4061 95
rect 4187 -196 4219 95
rect 4345 -196 4377 95
rect 4503 -196 4535 95
rect 4661 -196 4693 95
rect 4819 -196 4851 95
rect 4977 -196 5009 95
rect 5135 -196 5167 95
rect 5293 -196 5325 95
rect 5451 -196 5483 95
rect 5609 -196 5641 95
rect 5767 -196 5799 95
rect 5925 -196 5957 95
rect 6083 -196 6115 95
rect 6241 -196 6273 95
rect 6399 -196 6431 95
rect 6557 -196 6589 95
rect 3368 -233 6620 -196
rect 3368 -238 3534 -233
rect 3368 -300 3415 -238
rect 3368 -304 3534 -300
rect 3555 -304 3587 -233
rect 3713 -304 3745 -233
rect 3871 -304 3903 -233
rect 4029 -304 4061 -233
rect 4187 -304 4219 -233
rect 4345 -304 4377 -233
rect 4503 -304 4535 -233
rect 4661 -304 4693 -233
rect 4819 -304 4851 -233
rect 4977 -304 5009 -233
rect 5135 -304 5167 -233
rect 5293 -304 5325 -233
rect 5451 -304 5483 -233
rect 5609 -304 5641 -233
rect 5767 -304 5799 -233
rect 5925 -304 5957 -233
rect 6083 -304 6115 -233
rect 6241 -304 6273 -233
rect 6399 -304 6431 -233
rect 6557 -304 6589 -233
rect 3368 -341 6628 -304
rect 3368 -346 3534 -341
rect 3368 -628 3415 -346
rect 3368 -632 3534 -628
rect 3555 -632 3587 -341
rect 3713 -632 3745 -341
rect 3871 -632 3903 -341
rect 4029 -632 4061 -341
rect 4187 -632 4219 -341
rect 4345 -632 4377 -341
rect 4503 -632 4535 -341
rect 4661 -632 4693 -341
rect 4819 -632 4851 -341
rect 4977 -632 5009 -341
rect 5135 -632 5167 -341
rect 5293 -632 5325 -341
rect 5451 -632 5483 -341
rect 5609 -632 5641 -341
rect 5767 -632 5799 -341
rect 5925 -632 5957 -341
rect 6083 -632 6115 -341
rect 6241 -632 6273 -341
rect 6399 -632 6431 -341
rect 6557 -632 6589 -341
rect 3368 -669 6620 -632
rect 3368 -674 3534 -669
rect 3368 -736 3415 -674
rect 3368 -740 3534 -736
rect 3555 -740 3587 -669
rect 3713 -740 3745 -669
rect 3871 -740 3903 -669
rect 4029 -740 4061 -669
rect 4187 -740 4219 -669
rect 4345 -740 4377 -669
rect 4503 -740 4535 -669
rect 4661 -740 4693 -669
rect 4819 -740 4851 -669
rect 4977 -740 5009 -669
rect 5135 -740 5167 -669
rect 5293 -740 5325 -669
rect 5451 -740 5483 -669
rect 5609 -740 5641 -669
rect 5767 -740 5799 -669
rect 5925 -740 5957 -669
rect 6083 -740 6115 -669
rect 6241 -740 6273 -669
rect 6399 -740 6431 -669
rect 6557 -740 6589 -669
rect 3368 -777 6628 -740
rect 3368 -782 3534 -777
rect 3368 -1064 3415 -782
rect 3368 -1068 3534 -1064
rect 3555 -1068 3587 -777
rect 3713 -1068 3745 -777
rect 3871 -1068 3903 -777
rect 4029 -1068 4061 -777
rect 4187 -1068 4219 -777
rect 4345 -1068 4377 -777
rect 4503 -1068 4535 -777
rect 4661 -1068 4693 -777
rect 4819 -1068 4851 -777
rect 4977 -1068 5009 -777
rect 5135 -1068 5167 -777
rect 5293 -1068 5325 -777
rect 5451 -1068 5483 -777
rect 5609 -1068 5641 -777
rect 5767 -1068 5799 -777
rect 5925 -1068 5957 -777
rect 6083 -1068 6115 -777
rect 6241 -1068 6273 -777
rect 6399 -1068 6431 -777
rect 6557 -1068 6589 -777
rect 3368 -1105 6618 -1068
rect 3368 -1110 3534 -1105
rect 3713 -1110 3745 -1105
rect 3871 -1110 3903 -1105
rect 4029 -1110 4061 -1105
rect 4187 -1110 4219 -1105
rect 4345 -1110 4377 -1105
rect 4503 -1110 4535 -1105
rect 4661 -1110 4693 -1105
rect 4819 -1110 4851 -1105
rect 4977 -1110 5009 -1105
rect 5135 -1110 5167 -1105
rect 5293 -1110 5325 -1105
rect 5451 -1110 5483 -1105
rect 5609 -1110 5641 -1105
rect 5767 -1110 5799 -1105
rect 5925 -1110 5957 -1105
rect 6083 -1110 6115 -1105
rect 6241 -1110 6273 -1105
rect 6399 -1110 6431 -1105
rect 6557 -1110 6589 -1105
rect 3368 -1884 3415 -1110
rect 3462 -1188 6683 -1168
rect 3462 -1250 3502 -1188
rect 6650 -1200 6683 -1188
rect 6653 -1242 6683 -1200
rect 6650 -1250 6683 -1242
rect 3462 -1267 6683 -1250
rect 3555 -1346 3587 -1340
rect 3713 -1346 3745 -1340
rect 3871 -1346 3903 -1340
rect 4029 -1346 4061 -1340
rect 4187 -1346 4219 -1340
rect 4345 -1346 4377 -1340
rect 4503 -1346 4535 -1340
rect 4661 -1346 4693 -1340
rect 4819 -1346 4851 -1340
rect 4977 -1346 5009 -1340
rect 5135 -1346 5167 -1340
rect 5293 -1346 5325 -1340
rect 5451 -1346 5483 -1340
rect 5609 -1346 5641 -1340
rect 5767 -1346 5799 -1340
rect 5925 -1346 5957 -1340
rect 6083 -1346 6115 -1340
rect 6241 -1346 6273 -1340
rect 6399 -1346 6431 -1340
rect 6557 -1346 6589 -1340
rect 3517 -1383 6628 -1346
rect 3555 -1673 3587 -1383
rect 3713 -1673 3745 -1383
rect 3871 -1673 3903 -1383
rect 4029 -1673 4061 -1383
rect 4187 -1673 4219 -1383
rect 4345 -1673 4377 -1383
rect 4503 -1673 4535 -1383
rect 4661 -1673 4693 -1383
rect 4819 -1673 4851 -1383
rect 4977 -1673 5009 -1383
rect 5135 -1673 5167 -1383
rect 5293 -1673 5325 -1383
rect 5451 -1673 5483 -1383
rect 5609 -1673 5641 -1383
rect 5767 -1673 5799 -1383
rect 5925 -1673 5957 -1383
rect 6083 -1673 6115 -1383
rect 6241 -1673 6273 -1383
rect 6399 -1673 6431 -1383
rect 6557 -1673 6589 -1383
rect 3514 -1710 6625 -1673
rect 3555 -1714 3587 -1710
rect 3713 -1714 3745 -1710
rect 3871 -1714 3903 -1710
rect 4029 -1714 4061 -1710
rect 4187 -1714 4219 -1710
rect 4345 -1714 4377 -1710
rect 4503 -1714 4535 -1710
rect 4661 -1714 4693 -1710
rect 4819 -1714 4851 -1710
rect 4977 -1714 5009 -1710
rect 5135 -1714 5167 -1710
rect 5293 -1714 5325 -1710
rect 5451 -1714 5483 -1710
rect 5609 -1714 5641 -1710
rect 5767 -1714 5799 -1710
rect 3514 -1799 5822 -1784
rect 3514 -1834 3540 -1799
rect 5787 -1834 5822 -1799
rect 3514 -1848 5822 -1834
rect 3368 -1931 5021 -1884
rect 3309 -1975 4903 -1969
rect 3309 -2023 3338 -1975
rect 4871 -2023 4903 -1975
rect 3309 -2030 4903 -2023
rect 3309 -2255 3320 -2030
rect 4974 -2100 5021 -1931
rect 5066 -1974 5843 -1967
rect 5066 -2021 5095 -1974
rect 5809 -2021 5843 -1974
rect 5066 -2035 5843 -2021
rect 5878 -2100 5916 -1710
rect 5925 -1714 5957 -1710
rect 6083 -1714 6115 -1710
rect 6241 -1714 6273 -1710
rect 6399 -1714 6431 -1710
rect 6557 -1714 6589 -1710
rect 6773 -1785 6793 5004
rect 5956 -1801 6793 -1785
rect 5956 -1835 5977 -1801
rect 6669 -1835 6793 -1801
rect 5956 -1848 6793 -1835
rect 6773 -1968 6793 -1848
rect 5959 -1978 6793 -1968
rect 5959 -2025 5986 -1978
rect 6662 -2025 6793 -1978
rect 5959 -2035 6793 -2025
rect 4954 -2119 5042 -2100
rect 3213 -4457 3320 -2255
rect 3454 -2452 3491 -2205
rect 3550 -2452 3581 -2143
rect 3708 -2452 3739 -2143
rect 3866 -2452 3897 -2143
rect 3454 -2490 3937 -2452
rect 3365 -4239 3412 -3012
rect 3450 -3809 3490 -2916
rect 3549 -3550 3586 -2490
rect 4292 -2543 4323 -2141
rect 4450 -2543 4481 -2132
rect 3729 -2574 4481 -2543
rect 4450 -2732 4481 -2574
rect 4608 -2666 4639 -2128
rect 4766 -2666 4797 -2128
rect 4954 -2535 4970 -2119
rect 5029 -2535 5042 -2119
rect 5858 -2116 5935 -2100
rect 5192 -2449 5223 -2142
rect 5350 -2449 5381 -2142
rect 5508 -2449 5539 -2142
rect 5577 -2449 5628 -2406
rect 5666 -2449 5697 -2142
rect 5158 -2492 5736 -2449
rect 4954 -2551 5042 -2535
rect 5858 -2539 5869 -2116
rect 5924 -2539 5935 -2116
rect 6094 -2451 6125 -2136
rect 6252 -2451 6283 -2136
rect 6410 -2449 6441 -2136
rect 6481 -2449 6527 -2374
rect 6568 -2449 6599 -2136
rect 6379 -2451 6629 -2449
rect 6061 -2492 6633 -2451
rect 6379 -2495 6629 -2492
rect 6773 -2512 6793 -2035
rect 6832 -1142 6877 5063
rect 6950 -1142 6987 5187
rect 6832 -1260 6987 -1142
rect 6832 -1943 6877 -1260
rect 6950 -1943 6987 -1260
rect 6832 -2052 6987 -1943
rect 6832 -2512 6877 -2052
rect 6773 -2538 6877 -2512
rect 5858 -2553 5935 -2539
rect 6950 -2558 6987 -2052
rect 7030 -2558 7051 5187
rect 6950 -2585 7051 -2558
rect 6782 -2649 7016 -2641
rect 5863 -2666 5894 -2665
rect 6782 -2666 6791 -2649
rect 4608 -2697 6791 -2666
rect 4450 -2763 5657 -2732
rect 3674 -2981 3832 -2979
rect 3674 -3025 4261 -2981
rect 3674 -3026 3832 -3025
rect 3709 -3027 3832 -3026
rect 4109 -3027 4261 -3025
rect 3709 -3328 3740 -3027
rect 4139 -3330 4170 -3027
rect 4209 -3054 4261 -3027
rect 4568 -3329 4599 -2763
rect 4726 -2846 5041 -2815
rect 4726 -3295 4757 -2846
rect 5157 -3001 5188 -2987
rect 4709 -3332 4772 -3295
rect 3684 -3419 5119 -3398
rect 3684 -3470 3727 -3419
rect 5077 -3470 5119 -3419
rect 3684 -3489 5119 -3470
rect 5156 -3440 5191 -3001
rect 5626 -3326 5657 -2763
rect 5863 -2988 5894 -2697
rect 6782 -2715 6791 -2697
rect 7006 -2715 7016 -2649
rect 6782 -2723 7016 -2715
rect 6647 -2836 7020 -2809
rect 5863 -3327 5897 -2988
rect 5863 -3331 5894 -3327
rect 6336 -3440 6367 -2989
rect 6494 -3440 6525 -2989
rect 5156 -3475 6525 -3440
rect 6647 -3444 6687 -2836
rect 6742 -3444 7020 -2836
rect 3549 -3587 5731 -3550
rect 3541 -3636 5636 -3623
rect 3541 -3688 3588 -3636
rect 5602 -3640 5636 -3636
rect 5605 -3677 5636 -3640
rect 5602 -3688 5636 -3677
rect 3541 -3717 5636 -3688
rect 3541 -3724 3798 -3717
rect 3450 -3849 3668 -3809
rect 3615 -4359 3651 -4073
rect 3756 -4132 3798 -3724
rect 3755 -4197 3798 -4132
rect 3836 -3724 5636 -3717
rect 3836 -3730 4056 -3724
rect 3836 -4197 3973 -3730
rect 3755 -4198 3973 -4197
rect 4014 -4191 4056 -3730
rect 4225 -3823 4791 -3777
rect 4327 -3855 4373 -3823
rect 4643 -3855 4689 -3823
rect 4254 -4087 4285 -3864
rect 4412 -4087 4443 -3864
rect 4570 -4087 4601 -3864
rect 4728 -4087 4759 -3864
rect 4014 -4198 5103 -4191
rect 3755 -4221 5103 -4198
rect 3755 -4269 4160 -4221
rect 5053 -4269 5103 -4221
rect 3755 -4304 5103 -4269
rect 3755 -4437 4056 -4304
rect 5158 -4359 5189 -3785
rect 5262 -4333 5325 -3860
rect 5389 -4255 5517 -3854
rect 5588 -4124 5619 -3815
rect 5694 -4056 5731 -3587
rect 5803 -4015 5838 -3475
rect 6647 -3546 7020 -3444
rect 5956 -3563 7020 -3546
rect 5956 -3702 5984 -3563
rect 6676 -3653 7020 -3563
rect 6676 -3702 6688 -3653
rect 5956 -3726 6688 -3702
rect 6017 -4200 6048 -3784
rect 6175 -4200 6206 -3784
rect 6333 -4200 6364 -3784
rect 6491 -4101 6522 -3784
rect 6490 -4123 6522 -4101
rect 6490 -4200 6521 -4123
rect 6017 -4206 6521 -4200
rect 6017 -4231 6032 -4206
rect 6018 -4258 6032 -4231
rect 6497 -4231 6521 -4206
rect 6497 -4258 6506 -4231
rect 6018 -4268 6506 -4258
rect 6647 -4261 6688 -3726
rect 6743 -4261 7020 -3653
rect 6647 -4302 7020 -4261
rect 5262 -4396 6627 -4333
rect 3213 -4754 3223 -4457
rect 3310 -4754 3320 -4457
rect 3372 -4460 6232 -4437
rect 3372 -4523 3416 -4460
rect 6183 -4523 6232 -4460
rect 3372 -4545 6232 -4523
rect 3213 -4776 3320 -4754
rect 3293 -4898 3400 -4861
rect 3467 -4868 3899 -4632
rect 6300 -4676 6627 -4396
rect 6806 -4436 7020 -4302
rect 6806 -4457 6867 -4436
rect 3293 -5043 3322 -4898
rect 3369 -5043 3400 -4898
rect 3293 -5092 3400 -5043
rect 3451 -4973 3887 -4958
rect 3451 -5028 3468 -4973
rect 3871 -5028 3887 -4973
rect 3451 -5044 3887 -5028
rect 6200 -5034 6632 -4798
rect 6806 -5092 6823 -4457
rect 3246 -5116 6823 -5092
rect 3246 -5177 3269 -5116
rect 6803 -5121 6823 -5116
rect 6863 -5121 6867 -4457
rect 6803 -5132 6867 -5121
rect 6921 -5132 7020 -4436
rect 6803 -5177 7020 -5132
rect 3246 -5198 7020 -5177
rect 3042 -5359 3146 -5348
rect 3042 -5387 7058 -5359
rect 3042 -5441 3118 -5387
rect 6980 -5441 7058 -5387
rect 3042 -5471 7058 -5441
rect 7141 -5538 7164 5389
rect 2863 -5568 7164 -5538
rect 2863 -5614 3011 -5568
rect 7122 -5570 7164 -5568
rect 7210 -5570 7240 5438
rect 7122 -5614 7240 -5570
rect 2863 -5640 7240 -5614
<< via1 >>
rect 3407 5066 6621 5078
rect 3407 5031 6621 5066
rect 3407 5024 6621 5031
rect 3223 4770 3309 4788
rect 3223 -1823 3246 4770
rect 3246 -1823 3300 4770
rect 3300 -1823 3309 4770
rect 3223 -2255 3309 -1823
rect 3502 -1200 6650 -1188
rect 3502 -1242 3509 -1200
rect 3509 -1242 6650 -1200
rect 3502 -1250 6650 -1242
rect 4970 -2535 5029 -2119
rect 5869 -2539 5924 -2116
rect 6791 -2715 7006 -2649
rect 3588 -3640 5602 -3636
rect 3588 -3677 3597 -3640
rect 3597 -3677 5602 -3640
rect 3588 -3688 5602 -3677
rect 5984 -3702 6676 -3563
rect 6032 -4258 6497 -4206
rect 3223 -4754 3310 -4457
rect 3416 -4471 6183 -4460
rect 3416 -4507 3427 -4471
rect 3427 -4507 6153 -4471
rect 6153 -4507 6183 -4471
rect 3416 -4523 6183 -4507
rect 3468 -5028 3871 -4973
rect 3269 -5124 6803 -5116
rect 3269 -5161 3317 -5124
rect 3317 -5161 6782 -5124
rect 6782 -5161 6803 -5124
rect 6867 -5132 6921 -4436
rect 3269 -5177 6803 -5161
<< metal2 >>
rect 3120 5078 6663 5142
rect 3120 5024 3407 5078
rect 6621 5024 6663 5078
rect 3120 4984 6663 5024
rect 3120 4788 3412 4984
rect 6724 4939 7016 5142
rect 3459 4810 7016 4939
rect 3120 -2035 3223 4788
rect 3121 -2255 3223 -2035
rect 3309 4680 3412 4788
rect 3309 4551 6688 4680
rect 3309 4244 3412 4551
rect 6724 4503 7016 4810
rect 3459 4374 7016 4503
rect 3309 4115 6688 4244
rect 3309 3808 3412 4115
rect 6724 4067 7016 4374
rect 3459 3938 7016 4067
rect 3309 3679 6688 3808
rect 3309 3372 3412 3679
rect 6724 3631 7016 3938
rect 3459 3502 7016 3631
rect 3309 3243 6688 3372
rect 3309 2936 3412 3243
rect 6724 3195 7016 3502
rect 3459 3066 7016 3195
rect 3309 2807 6688 2936
rect 3309 2500 3412 2807
rect 6724 2759 7016 3066
rect 3459 2630 7016 2759
rect 3309 2371 6688 2500
rect 3309 2064 3412 2371
rect 6724 2323 7016 2630
rect 3459 2194 7016 2323
rect 3309 1935 6688 2064
rect 3309 1628 3412 1935
rect 6724 1887 7016 2194
rect 3459 1758 7016 1887
rect 3309 1499 6688 1628
rect 3309 1192 3412 1499
rect 6724 1451 7016 1758
rect 3459 1322 7016 1451
rect 3309 1063 6688 1192
rect 3309 756 3412 1063
rect 6724 1015 7016 1322
rect 3459 886 7016 1015
rect 3309 627 6688 756
rect 3309 320 3412 627
rect 6724 579 7016 886
rect 3459 450 7016 579
rect 3309 191 6688 320
rect 3309 -116 3412 191
rect 6724 143 7016 450
rect 3459 14 7016 143
rect 3309 -245 6688 -116
rect 3309 -552 3412 -245
rect 6724 -293 7016 14
rect 3459 -422 7016 -293
rect 3309 -681 6688 -552
rect 3309 -988 3412 -681
rect 6724 -729 7016 -422
rect 3459 -858 7016 -729
rect 3309 -1117 6688 -988
rect 3309 -1165 3412 -1117
rect 3309 -1188 6686 -1165
rect 3309 -1250 3502 -1188
rect 6650 -1250 6686 -1188
rect 3309 -1271 6686 -1250
rect 3309 -1592 3412 -1271
rect 6724 -1333 7016 -858
rect 3462 -1462 7016 -1333
rect 3309 -1721 6691 -1592
rect 3309 -1785 3412 -1721
rect 6724 -1765 7016 -1462
rect 3309 -1862 6692 -1785
rect 3309 -2035 6691 -1862
rect 3309 -2177 3412 -2035
rect 4954 -2119 5042 -2100
rect 3309 -2178 3421 -2177
rect 3309 -2255 4011 -2178
rect 3121 -2265 4011 -2255
rect 4068 -2264 4906 -2180
rect 4068 -2351 4152 -2264
rect 3436 -2435 4152 -2351
rect 3120 -2530 3320 -2460
rect 4356 -2528 4419 -2292
rect 3120 -2592 3727 -2530
rect 3964 -2591 4419 -2528
rect 3120 -2660 3320 -2592
rect 3446 -2804 3489 -2592
rect 3964 -2780 4027 -2591
rect 4665 -2653 4728 -2292
rect 4954 -2531 4970 -2119
rect 3773 -2843 4027 -2780
rect 4203 -2716 4728 -2653
rect 4867 -2535 4970 -2531
rect 5029 -2531 5042 -2119
rect 5073 -2178 5158 -2035
rect 5858 -2116 5935 -2100
rect 5073 -2263 5797 -2178
rect 5255 -2531 5321 -2292
rect 5029 -2535 5321 -2531
rect 4867 -2597 5321 -2535
rect 3773 -2979 3836 -2843
rect 3389 -3044 3836 -2979
rect 3592 -3381 3704 -3114
rect 3773 -3180 3836 -3044
rect 4014 -3381 4126 -3113
rect 4203 -3182 4266 -2716
rect 4867 -2764 4933 -2597
rect 5570 -2684 5636 -2291
rect 5858 -2533 5869 -2116
rect 4472 -2830 4933 -2764
rect 5022 -2812 5076 -2684
rect 5185 -2750 5636 -2684
rect 5775 -2539 5869 -2533
rect 5924 -2533 5935 -2116
rect 5973 -2178 6058 -2035
rect 5973 -2263 6697 -2178
rect 5973 -2264 6060 -2263
rect 5996 -2323 6002 -2264
rect 6054 -2323 6060 -2264
rect 6155 -2533 6221 -2292
rect 6312 -2323 6318 -2263
rect 6370 -2323 6376 -2263
rect 5924 -2539 6221 -2533
rect 5775 -2599 6221 -2539
rect 4472 -3184 4538 -2830
rect 5185 -2898 5251 -2750
rect 4793 -2964 5251 -2898
rect 4605 -3227 4717 -3114
rect 4793 -3186 4859 -2964
rect 5775 -3008 5841 -2599
rect 6470 -2693 6536 -2291
rect 6629 -2323 6635 -2263
rect 6687 -2323 6693 -2263
rect 5484 -3074 5841 -3008
rect 5968 -2759 6536 -2693
rect 6782 -2649 7016 -1765
rect 6782 -2715 6791 -2649
rect 7006 -2715 7016 -2649
rect 4605 -3317 5127 -3227
rect 5206 -3381 5309 -3126
rect 5484 -3178 5550 -3074
rect 5708 -3227 5820 -3113
rect 5968 -3180 6034 -2759
rect 6101 -3083 6611 -2993
rect 6101 -3227 6191 -3083
rect 5708 -3317 6191 -3227
rect 6377 -3381 6480 -3127
rect 3122 -3563 6695 -3381
rect 3122 -3636 5984 -3563
rect 3122 -3688 3588 -3636
rect 5602 -3688 5984 -3636
rect 3122 -3702 5984 -3688
rect 6676 -3702 6695 -3563
rect 3122 -3899 6695 -3702
rect 6782 -4017 7016 -2715
rect 4091 -4130 5863 -4017
rect 5941 -4130 7016 -4017
rect 3124 -4357 3324 -4193
rect 3414 -4206 6512 -4195
rect 3414 -4239 6032 -4206
rect 6011 -4258 6032 -4239
rect 6497 -4239 6512 -4206
rect 6497 -4258 6511 -4239
rect 6011 -4259 6511 -4258
rect 3124 -4393 5189 -4357
rect 6806 -4436 7020 -4356
rect 6806 -4437 6867 -4436
rect 3213 -4457 3320 -4437
rect 3213 -4754 3223 -4457
rect 3310 -4754 3320 -4457
rect 3372 -4460 6867 -4437
rect 3372 -4523 3416 -4460
rect 6183 -4523 6867 -4460
rect 3372 -4545 6867 -4523
rect 3213 -4958 3320 -4754
rect 3213 -4973 3887 -4958
rect 3213 -5028 3468 -4973
rect 3871 -5028 3887 -4973
rect 3213 -5042 3887 -5028
rect 6806 -5092 6867 -4545
rect 3246 -5116 6867 -5092
rect 3246 -5177 3269 -5116
rect 6803 -5132 6867 -5116
rect 6921 -5132 7020 -4436
rect 6803 -5177 7020 -5132
rect 3246 -5198 7020 -5177
use amp_via_2cut  amp_via_2cut_0
timestamp 1717613630
transform 0 1 11393 -1 0 15277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_1
timestamp 1717613630
transform 0 1 11551 -1 0 15189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_2
timestamp 1717613630
transform 0 1 11867 -1 0 15189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_3
timestamp 1717613630
transform 0 1 11709 -1 0 15277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_4
timestamp 1717613630
transform 0 1 13447 -1 0 14584
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_5
timestamp 1717613630
transform 0 1 13289 -1 0 14672
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_6
timestamp 1717613630
transform 0 1 12183 -1 0 14584
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_7
timestamp 1717613630
transform 0 1 12025 -1 0 14672
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_8
timestamp 1717613630
transform 0 1 12499 -1 0 14584
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_9
timestamp 1717613630
transform 0 1 12341 -1 0 14672
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_10
timestamp 1717613630
transform 0 1 12815 -1 0 14584
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_11
timestamp 1717613630
transform 0 1 12657 -1 0 14672
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_12
timestamp 1717613630
transform 0 1 13131 -1 0 14584
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_13
timestamp 1717613630
transform 0 1 12973 -1 0 14672
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_14
timestamp 1717613630
transform 0 1 14395 -1 0 15189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_15
timestamp 1717613630
transform 0 1 14553 -1 0 15277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_16
timestamp 1717613630
transform 0 1 13763 -1 0 15189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_17
timestamp 1717613630
transform 0 1 13605 -1 0 15277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_18
timestamp 1717613630
transform 0 1 14079 -1 0 15189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_19
timestamp 1717613630
transform 0 1 13921 -1 0 15277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_20
timestamp 1717613630
transform 0 1 14237 -1 0 15277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_21
timestamp 1717613630
transform 0 1 11867 -1 0 14584
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_22
timestamp 1717613630
transform 0 1 11709 -1 0 14672
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_23
timestamp 1717613630
transform 0 1 11393 -1 0 14672
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_24
timestamp 1717613630
transform 0 1 11862 1 0 -18417
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_25
timestamp 1717613630
transform 0 1 12341 -1 0 15277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_26
timestamp 1717613630
transform 0 1 12025 -1 0 15277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_27
timestamp 1717613630
transform 0 1 12183 -1 0 15189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_28
timestamp 1717613630
transform 0 1 12657 -1 0 15277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_29
timestamp 1717613630
transform 0 1 12815 -1 0 15189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_30
timestamp 1717613630
transform 0 1 12499 -1 0 15189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_31
timestamp 1717613630
transform 0 1 13289 -1 0 15277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_32
timestamp 1717613630
transform 0 1 13131 -1 0 15189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_33
timestamp 1717613630
transform 0 1 12973 -1 0 15277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_34
timestamp 1717613630
transform 0 1 13447 -1 0 15189
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_35
timestamp 1717613630
transform 0 1 14553 -1 0 14672
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_36
timestamp 1717613630
transform 0 1 14395 -1 0 14584
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_37
timestamp 1717613630
transform 0 1 14237 -1 0 14672
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_38
timestamp 1717613630
transform 0 1 14079 -1 0 14584
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_39
timestamp 1717613630
transform 0 1 13921 -1 0 14672
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_40
timestamp 1717613630
transform 0 1 13763 -1 0 14584
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_41
timestamp 1717613630
transform 0 1 13605 -1 0 14672
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_42
timestamp 1717613630
transform 0 1 11709 -1 0 15713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_43
timestamp 1717613630
transform 0 1 11867 -1 0 15625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_44
timestamp 1717613630
transform 0 1 11393 -1 0 15713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_45
timestamp 1717613630
transform 0 1 11551 -1 0 15625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_46
timestamp 1717613630
transform 0 1 13447 -1 0 15625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_47
timestamp 1717613630
transform 0 1 13289 -1 0 15713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_48
timestamp 1717613630
transform 0 1 13131 -1 0 15625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_49
timestamp 1717613630
transform 0 1 12973 -1 0 15713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_50
timestamp 1717613630
transform 0 1 12657 -1 0 15713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_51
timestamp 1717613630
transform 0 1 12815 -1 0 15625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_52
timestamp 1717613630
transform 0 1 12341 -1 0 15713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_53
timestamp 1717613630
transform 0 1 12499 -1 0 15625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_54
timestamp 1717613630
transform 0 1 12025 -1 0 15713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_55
timestamp 1717613630
transform 0 1 12183 -1 0 15625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_56
timestamp 1717613630
transform 0 1 14553 -1 0 15713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_57
timestamp 1717613630
transform 0 1 14395 -1 0 15625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_58
timestamp 1717613630
transform 0 1 14237 -1 0 15713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_59
timestamp 1717613630
transform 0 1 14079 -1 0 15625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_60
timestamp 1717613630
transform 0 1 13921 -1 0 15713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_61
timestamp 1717613630
transform 0 1 13763 -1 0 15625
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_62
timestamp 1717613630
transform 0 1 13605 -1 0 15713
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_63
timestamp 1717613630
transform 0 1 14553 -1 0 17021
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_64
timestamp 1717613630
transform 0 1 14395 -1 0 16933
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_65
timestamp 1717613630
transform 0 1 14237 -1 0 17021
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_66
timestamp 1717613630
transform 0 1 14079 -1 0 16933
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_67
timestamp 1717613630
transform 0 1 13921 -1 0 17021
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_68
timestamp 1717613630
transform 0 1 13763 -1 0 16933
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_69
timestamp 1717613630
transform 0 1 13605 -1 0 17021
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_70
timestamp 1717613630
transform 0 1 13447 -1 0 16933
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_71
timestamp 1717613630
transform 0 1 13289 -1 0 16585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_72
timestamp 1717613630
transform 0 1 13131 -1 0 16497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_73
timestamp 1717613630
transform 0 1 12973 -1 0 16585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_74
timestamp 1717613630
transform 0 1 12657 -1 0 16585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_75
timestamp 1717613630
transform 0 1 12815 -1 0 16497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_76
timestamp 1717613630
transform 0 1 12341 -1 0 16585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_77
timestamp 1717613630
transform 0 1 12499 -1 0 16497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_78
timestamp 1717613630
transform 0 1 12025 -1 0 16585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_79
timestamp 1717613630
transform 0 1 12183 -1 0 16497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_80
timestamp 1717613630
transform 0 1 11709 -1 0 17021
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_81
timestamp 1717613630
transform 0 1 11867 -1 0 16933
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_82
timestamp 1717613630
transform 0 1 11393 -1 0 17021
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_83
timestamp 1717613630
transform 0 1 11551 -1 0 16933
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_84
timestamp 1717613630
transform 0 1 11551 -1 0 16061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_85
timestamp 1717613630
transform 0 1 11393 -1 0 16149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_86
timestamp 1717613630
transform 0 1 11867 -1 0 16061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_87
timestamp 1717613630
transform 0 1 11709 -1 0 16149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_88
timestamp 1717613630
transform 0 1 12183 -1 0 16061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_89
timestamp 1717613630
transform 0 1 12025 -1 0 16149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_90
timestamp 1717613630
transform 0 1 12499 -1 0 16061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_91
timestamp 1717613630
transform 0 1 12341 -1 0 16149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_92
timestamp 1717613630
transform 0 1 12815 -1 0 16061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_93
timestamp 1717613630
transform 0 1 12657 -1 0 16149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_94
timestamp 1717613630
transform 0 1 12973 -1 0 16149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_95
timestamp 1717613630
transform 0 1 13131 -1 0 16061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_96
timestamp 1717613630
transform 0 1 13289 -1 0 16149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_97
timestamp 1717613630
transform 0 1 13447 -1 0 16061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_98
timestamp 1717613630
transform 0 1 13605 -1 0 16149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_99
timestamp 1717613630
transform 0 1 13763 -1 0 16061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_100
timestamp 1717613630
transform 0 1 13921 -1 0 16149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_101
timestamp 1717613630
transform 0 1 14079 -1 0 16061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_102
timestamp 1717613630
transform 0 1 14237 -1 0 16149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_103
timestamp 1717613630
transform 0 1 14395 -1 0 16061
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_104
timestamp 1717613630
transform 0 1 14553 -1 0 16149
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_105
timestamp 1717613630
transform 0 1 11709 -1 0 16585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_106
timestamp 1717613630
transform 0 1 11867 -1 0 16497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_107
timestamp 1717613630
transform 0 1 11393 -1 0 16585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_108
timestamp 1717613630
transform 0 1 11551 -1 0 16497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_109
timestamp 1717613630
transform 0 1 12183 -1 0 16933
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_110
timestamp 1717613630
transform 0 1 12499 -1 0 16933
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_111
timestamp 1717613630
transform 0 1 12815 -1 0 16933
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_112
timestamp 1717613630
transform 0 1 13131 -1 0 16933
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_113
timestamp 1717613630
transform 0 1 12025 -1 0 17021
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_114
timestamp 1717613630
transform 0 1 12341 -1 0 17021
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_115
timestamp 1717613630
transform 0 1 12657 -1 0 17021
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_116
timestamp 1717613630
transform 0 1 13289 -1 0 17021
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_117
timestamp 1717613630
transform 0 1 12973 -1 0 17021
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_118
timestamp 1717613630
transform 0 1 14553 -1 0 16585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_119
timestamp 1717613630
transform 0 1 14395 -1 0 16497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_120
timestamp 1717613630
transform 0 1 14237 -1 0 16585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_121
timestamp 1717613630
transform 0 1 14079 -1 0 16497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_122
timestamp 1717613630
transform 0 1 13921 -1 0 16585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_123
timestamp 1717613630
transform 0 1 13763 -1 0 16497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_124
timestamp 1717613630
transform 0 1 13605 -1 0 16585
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_125
timestamp 1717613630
transform 0 1 13447 -1 0 16497
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_126
timestamp 1717613630
transform 0 1 11551 -1 0 17369
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_127
timestamp 1717613630
transform 0 1 11867 -1 0 17369
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_128
timestamp 1717613630
transform 0 1 12183 -1 0 17369
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_129
timestamp 1717613630
transform 0 1 12499 -1 0 17369
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_130
timestamp 1717613630
transform 0 1 12815 -1 0 17369
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_131
timestamp 1717613630
transform 0 1 13131 -1 0 17369
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_132
timestamp 1717613630
transform 0 1 13447 -1 0 17369
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_133
timestamp 1717613630
transform 0 1 13763 -1 0 17369
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_134
timestamp 1717613630
transform 0 1 14079 -1 0 17369
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_135
timestamp 1717613630
transform 0 1 14395 -1 0 17369
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_136
timestamp 1717613630
transform 0 1 11709 -1 0 18329
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_137
timestamp 1717613630
transform 0 1 11393 -1 0 18329
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_138
timestamp 1717613630
transform 0 1 13289 -1 0 17893
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_139
timestamp 1717613630
transform 0 1 12973 -1 0 17893
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_140
timestamp 1717613630
transform 0 1 12657 -1 0 17893
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_141
timestamp 1717613630
transform 0 1 12341 -1 0 17893
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_142
timestamp 1717613630
transform 0 1 12025 -1 0 17893
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_143
timestamp 1717613630
transform 0 1 14553 -1 0 18329
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_144
timestamp 1717613630
transform 0 1 14237 -1 0 18329
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_145
timestamp 1717613630
transform 0 1 13921 -1 0 18329
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_146
timestamp 1717613630
transform 0 1 13605 -1 0 18329
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_147
timestamp 1717613630
transform 0 1 11867 -1 0 18241
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_148
timestamp 1717613630
transform 0 1 11551 -1 0 18241
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_149
timestamp 1717613630
transform 0 1 11709 -1 0 17457
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_150
timestamp 1717613630
transform 0 1 11393 -1 0 17457
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_151
timestamp 1717613630
transform 0 1 13131 -1 0 17805
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_152
timestamp 1717613630
transform 0 1 12815 -1 0 17805
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_153
timestamp 1717613630
transform 0 1 12499 -1 0 17805
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_154
timestamp 1717613630
transform 0 1 12183 -1 0 17805
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_155
timestamp 1717613630
transform 0 1 13289 -1 0 17457
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_156
timestamp 1717613630
transform 0 1 12973 -1 0 17457
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_157
timestamp 1717613630
transform 0 1 12657 -1 0 17457
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_158
timestamp 1717613630
transform 0 1 12341 -1 0 17457
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_159
timestamp 1717613630
transform 0 1 12025 -1 0 17457
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_160
timestamp 1717613630
transform 0 1 14395 -1 0 18241
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_161
timestamp 1717613630
transform 0 1 14079 -1 0 18241
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_162
timestamp 1717613630
transform 0 1 13763 -1 0 18241
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_163
timestamp 1717613630
transform 0 1 13447 -1 0 18241
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_164
timestamp 1717613630
transform 0 1 14553 -1 0 17457
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_165
timestamp 1717613630
transform 0 1 14237 -1 0 17457
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_166
timestamp 1717613630
transform 0 1 13921 -1 0 17457
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_167
timestamp 1717613630
transform 0 1 13605 -1 0 17457
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_168
timestamp 1717613630
transform 0 1 11709 -1 0 17893
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_169
timestamp 1717613630
transform 0 1 11867 -1 0 17805
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_170
timestamp 1717613630
transform 0 1 11393 -1 0 17893
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_171
timestamp 1717613630
transform 0 1 11551 -1 0 17805
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_172
timestamp 1717613630
transform 0 1 12025 -1 0 18329
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_173
timestamp 1717613630
transform 0 1 12183 -1 0 18241
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_174
timestamp 1717613630
transform 0 1 12657 -1 0 18329
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_175
timestamp 1717613630
transform 0 1 12341 -1 0 18329
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_176
timestamp 1717613630
transform 0 1 12499 -1 0 18241
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_177
timestamp 1717613630
transform 0 1 12973 -1 0 18329
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_178
timestamp 1717613630
transform 0 1 12815 -1 0 18241
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_179
timestamp 1717613630
transform 0 1 13289 -1 0 18329
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_180
timestamp 1717613630
transform 0 1 13131 -1 0 18241
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_181
timestamp 1717613630
transform 0 1 14553 -1 0 17893
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_182
timestamp 1717613630
transform 0 1 14395 -1 0 17805
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_183
timestamp 1717613630
transform 0 1 14237 -1 0 17893
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_184
timestamp 1717613630
transform 0 1 14079 -1 0 17805
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_185
timestamp 1717613630
transform 0 1 13921 -1 0 17893
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_186
timestamp 1717613630
transform 0 1 13763 -1 0 17805
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_187
timestamp 1717613630
transform 0 1 13605 -1 0 17893
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_188
timestamp 1717613630
transform 0 1 13447 -1 0 17805
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_189
timestamp 1717613630
transform 0 1 11867 -1 0 18677
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_190
timestamp 1717613630
transform 0 1 11551 -1 0 18677
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_191
timestamp 1717613630
transform 0 1 11393 -1 0 18765
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_192
timestamp 1717613630
transform 0 1 11709 -1 0 18765
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_193
timestamp 1717613630
transform 0 1 12025 -1 0 18765
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_194
timestamp 1717613630
transform 0 1 12183 -1 0 18677
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_195
timestamp 1717613630
transform 0 1 12657 -1 0 18765
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_196
timestamp 1717613630
transform 0 1 12341 -1 0 18765
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_197
timestamp 1717613630
transform 0 1 12499 -1 0 18677
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_198
timestamp 1717613630
transform 0 1 12973 -1 0 18765
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_199
timestamp 1717613630
transform 0 1 12815 -1 0 18677
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_200
timestamp 1717613630
transform 0 1 13289 -1 0 18765
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_201
timestamp 1717613630
transform 0 1 13131 -1 0 18677
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_202
timestamp 1717613630
transform 0 1 13605 -1 0 18765
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_203
timestamp 1717613630
transform 0 1 13447 -1 0 18677
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_204
timestamp 1717613630
transform 0 1 13921 -1 0 18765
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_205
timestamp 1717613630
transform 0 1 13763 -1 0 18677
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_206
timestamp 1717613630
transform 0 1 14237 -1 0 18765
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_207
timestamp 1717613630
transform 0 1 14079 -1 0 18677
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_208
timestamp 1717613630
transform 0 1 14553 -1 0 18765
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_209
timestamp 1717613630
transform 0 1 14395 -1 0 18677
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_210
timestamp 1717613630
transform 0 1 11709 -1 0 20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_211
timestamp 1717613630
transform 0 1 11867 -1 0 19985
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_212
timestamp 1717613630
transform 0 1 11393 -1 0 20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_213
timestamp 1717613630
transform 0 1 11551 -1 0 19985
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_214
timestamp 1717613630
transform 0 1 13289 -1 0 19637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_215
timestamp 1717613630
transform 0 1 13131 -1 0 19549
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_216
timestamp 1717613630
transform 0 1 12973 -1 0 19637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_217
timestamp 1717613630
transform 0 1 12657 -1 0 19637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_218
timestamp 1717613630
transform 0 1 12815 -1 0 19549
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_219
timestamp 1717613630
transform 0 1 12341 -1 0 19637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_220
timestamp 1717613630
transform 0 1 12499 -1 0 19549
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_221
timestamp 1717613630
transform 0 1 12025 -1 0 19637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_222
timestamp 1717613630
transform 0 1 12183 -1 0 19549
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_223
timestamp 1717613630
transform 0 1 14553 -1 0 20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_224
timestamp 1717613630
transform 0 1 14395 -1 0 19985
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_225
timestamp 1717613630
transform 0 1 14237 -1 0 20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_226
timestamp 1717613630
transform 0 1 14079 -1 0 19985
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_227
timestamp 1717613630
transform 0 1 13921 -1 0 20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_228
timestamp 1717613630
transform 0 1 13763 -1 0 19985
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_229
timestamp 1717613630
transform 0 1 13605 -1 0 20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_230
timestamp 1717613630
transform 0 1 13447 -1 0 19985
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_231
timestamp 1717613630
transform 0 1 11709 -1 0 19201
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_232
timestamp 1717613630
transform 0 1 11867 -1 0 19113
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_233
timestamp 1717613630
transform 0 1 11393 -1 0 19201
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_234
timestamp 1717613630
transform 0 1 11551 -1 0 19113
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_235
timestamp 1717613630
transform 0 1 13289 -1 0 19201
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_236
timestamp 1717613630
transform 0 1 13131 -1 0 19113
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_237
timestamp 1717613630
transform 0 1 12973 -1 0 19201
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_238
timestamp 1717613630
transform 0 1 12657 -1 0 19201
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_239
timestamp 1717613630
transform 0 1 12815 -1 0 19113
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_240
timestamp 1717613630
transform 0 1 12341 -1 0 19201
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_241
timestamp 1717613630
transform 0 1 12499 -1 0 19113
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_242
timestamp 1717613630
transform 0 1 12025 -1 0 19201
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_243
timestamp 1717613630
transform 0 1 12183 -1 0 19113
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_244
timestamp 1717613630
transform 0 1 14553 -1 0 19201
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_245
timestamp 1717613630
transform 0 1 14395 -1 0 19113
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_246
timestamp 1717613630
transform 0 1 14237 -1 0 19201
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_247
timestamp 1717613630
transform 0 1 14079 -1 0 19113
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_248
timestamp 1717613630
transform 0 1 13921 -1 0 19201
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_249
timestamp 1717613630
transform 0 1 13763 -1 0 19113
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_250
timestamp 1717613630
transform 0 1 13605 -1 0 19201
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_251
timestamp 1717613630
transform 0 1 13447 -1 0 19113
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_252
timestamp 1717613630
transform 0 1 11709 -1 0 19637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_253
timestamp 1717613630
transform 0 1 11867 -1 0 19549
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_254
timestamp 1717613630
transform 0 1 11393 -1 0 19637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_255
timestamp 1717613630
transform 0 1 11551 -1 0 19549
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_256
timestamp 1717613630
transform 0 1 12025 -1 0 20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_257
timestamp 1717613630
transform 0 1 12183 -1 0 19985
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_258
timestamp 1717613630
transform 0 1 12341 -1 0 20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_259
timestamp 1717613630
transform 0 1 12499 -1 0 19985
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_260
timestamp 1717613630
transform 0 1 12657 -1 0 20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_261
timestamp 1717613630
transform 0 1 12815 -1 0 19985
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_262
timestamp 1717613630
transform 0 1 13289 -1 0 20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_263
timestamp 1717613630
transform 0 1 13131 -1 0 19985
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_264
timestamp 1717613630
transform 0 1 12973 -1 0 20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_265
timestamp 1717613630
transform 0 1 14553 -1 0 19637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_266
timestamp 1717613630
transform 0 1 14395 -1 0 19549
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_267
timestamp 1717613630
transform 0 1 14237 -1 0 19637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_268
timestamp 1717613630
transform 0 1 14079 -1 0 19549
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_269
timestamp 1717613630
transform 0 1 13921 -1 0 19637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_270
timestamp 1717613630
transform 0 1 13763 -1 0 19549
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_271
timestamp 1717613630
transform 0 1 13605 -1 0 19637
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_272
timestamp 1717613630
transform 0 1 13447 -1 0 19549
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_273
timestamp 1717613630
transform 0 1 11709 -1 0 20945
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_274
timestamp 1717613630
transform 0 1 11867 -1 0 20857
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_275
timestamp 1717613630
transform 0 1 11393 -1 0 20945
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_276
timestamp 1717613630
transform 0 1 11551 -1 0 20857
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_277
timestamp 1717613630
transform 0 1 13289 -1 0 20945
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_278
timestamp 1717613630
transform 0 1 13131 -1 0 20857
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_279
timestamp 1717613630
transform 0 1 12973 -1 0 20945
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_280
timestamp 1717613630
transform 0 1 12657 -1 0 20945
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_281
timestamp 1717613630
transform 0 1 12815 -1 0 20857
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_282
timestamp 1717613630
transform 0 1 12341 -1 0 20945
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_283
timestamp 1717613630
transform 0 1 12499 -1 0 20857
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_284
timestamp 1717613630
transform 0 1 12025 -1 0 20945
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_285
timestamp 1717613630
transform 0 1 12183 -1 0 20857
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_286
timestamp 1717613630
transform 0 1 14553 -1 0 20945
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_287
timestamp 1717613630
transform 0 1 14395 -1 0 20857
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_288
timestamp 1717613630
transform 0 1 14237 -1 0 20945
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_289
timestamp 1717613630
transform 0 1 14079 -1 0 20857
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_290
timestamp 1717613630
transform 0 1 13921 -1 0 20945
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_291
timestamp 1717613630
transform 0 1 13763 -1 0 20857
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_292
timestamp 1717613630
transform 0 1 13605 -1 0 20945
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_293
timestamp 1717613630
transform 0 1 13447 -1 0 20857
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_294
timestamp 1717613630
transform 0 1 11709 -1 0 20509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_295
timestamp 1717613630
transform 0 1 11867 -1 0 20421
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_296
timestamp 1717613630
transform 0 1 11393 -1 0 20509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_297
timestamp 1717613630
transform 0 1 11551 -1 0 20421
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_298
timestamp 1717613630
transform 0 1 13289 -1 0 20509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_299
timestamp 1717613630
transform 0 1 13131 -1 0 20421
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_300
timestamp 1717613630
transform 0 1 12973 -1 0 20509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_301
timestamp 1717613630
transform 0 1 12657 -1 0 20509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_302
timestamp 1717613630
transform 0 1 12815 -1 0 20421
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_303
timestamp 1717613630
transform 0 1 12341 -1 0 20509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_304
timestamp 1717613630
transform 0 1 12499 -1 0 20421
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_305
timestamp 1717613630
transform 0 1 12025 -1 0 20509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_306
timestamp 1717613630
transform 0 1 12183 -1 0 20421
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_307
timestamp 1717613630
transform 0 1 14553 -1 0 20509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_308
timestamp 1717613630
transform 0 1 14395 -1 0 20421
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_309
timestamp 1717613630
transform 0 1 14237 -1 0 20509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_310
timestamp 1717613630
transform 0 1 14079 -1 0 20421
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_311
timestamp 1717613630
transform 0 1 13921 -1 0 20509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_312
timestamp 1717613630
transform 0 1 13763 -1 0 20421
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_313
timestamp 1717613630
transform 0 1 13605 -1 0 20509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_314
timestamp 1717613630
transform 0 1 13447 -1 0 20421
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_315
timestamp 1717613630
transform 0 1 11551 -1 0 14584
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_316
timestamp 1717613630
transform 0 1 11705 1 0 -18509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_317
timestamp 1717613630
transform 0 1 11546 1 0 -18417
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_318
timestamp 1717613630
transform 0 1 12600 1 0 -18509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_319
timestamp 1717613630
transform 0 1 11975 1 0 -19352
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_320
timestamp 1717613630
transform 0 1 12445 1 0 -18417
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_321
timestamp 1717613630
transform 0 1 12129 1 0 -18417
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_322
timestamp 1717613630
transform 0 1 12762 1 0 -18417
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_323
timestamp 1717613630
transform 0 -1 -4514 -1 0 13121
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_324
timestamp 1717613630
transform 0 1 13417 1 0 -19274
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_325
timestamp 1717613630
transform 0 1 11705 1 0 -19278
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_326
timestamp 1717613630
transform 0 1 11546 1 0 -19351
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_327
timestamp 1717613630
transform 0 1 13189 1 0 -18508
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_328
timestamp 1717613630
transform 1 0 -12399 0 -1 -10463
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_329
timestamp 1717613630
transform 0 1 13344 1 0 -18417
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_330
timestamp 1717613630
transform 0 1 13028 1 0 -18417
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_331
timestamp 1717613630
transform 0 1 13661 1 0 -18417
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_332
timestamp 1717613630
transform 0 1 12287 1 0 -18508
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_333
timestamp 1717613630
transform 0 1 14402 1 0 -18509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_334
timestamp 1717613630
transform 0 1 14089 1 0 -18508
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_335
timestamp 1717613630
transform 0 1 13502 1 0 -18509
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_336
timestamp 1717613630
transform 0 1 14244 1 0 -18417
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_337
timestamp 1717613630
transform 0 1 13928 1 0 -18417
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_338
timestamp 1717613630
transform 0 1 14561 1 0 -18417
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_339
timestamp 1717613630
transform 0 1 12135 1 0 -19276
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_340
timestamp 1717613630
transform 0 1 12996 1 0 -20143
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_341
timestamp 1717613630
transform 0 1 12725 1 0 -19276
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_342
timestamp 1717613630
transform 0 1 13900 1 0 -19277
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_343
timestamp 1717613630
transform 0 1 13152 1 0 -19350
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_344
timestamp 1717613630
transform 0 1 13662 1 0 -19351
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_345
timestamp 1717613630
transform 0 1 12404 1 0 -19276
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_346
timestamp 1717613630
transform 0 1 12724 1 0 -20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_347
timestamp 1717613630
transform 0 1 12408 1 0 -20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_348
timestamp 1717613630
transform 0 1 12092 1 0 -20073
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_349
timestamp 1717613630
transform 0 1 12251 1 0 -20147
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_350
timestamp 1717613630
transform 1 0 -12728 0 -1 -12113
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_351
timestamp 1717613630
transform 0 1 13723 1 0 -20224
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_352
timestamp 1717613630
transform 1 0 -11107 0 -1 -10575
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_353
timestamp 1717613630
transform 1 0 -11104 0 -1 -10726
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_354
timestamp 1717613630
transform 0 1 12565 1 0 -19351
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_355
timestamp 1717613630
transform 0 1 14170 1 0 -19278
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_356
timestamp 1717613630
transform 0 1 12995 1 0 -19350
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_357
timestamp 1717613630
transform 0 1 14486 1 0 -19278
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_358
timestamp 1717613630
transform 0 1 14331 1 0 -19347
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_359
timestamp 1717613630
transform 1 0 -10520 0 -1 -12031
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_360
timestamp 1717613630
transform 1 0 -10993 0 -1 -12272
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_361
timestamp 1717613630
transform 0 1 13856 1 0 -20074
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_362
timestamp 1717613630
transform 0 1 14015 1 0 -20148
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_363
timestamp 1717613630
transform 0 1 14172 1 0 -20074
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_364
timestamp 1717613630
transform 0 1 14330 1 0 -20148
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_365
timestamp 1717613630
transform 0 1 14488 1 0 -20074
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_366
timestamp 1717613630
transform 0 1 12566 1 0 -20147
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_367
timestamp 1717613630
transform 1 0 -12513 0 -1 -12272
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_368
timestamp 1717613630
transform 0 -1 -4432 -1 0 13301
box 16088 -7932 16222 -7868
use amp_via_2cut  amp_via_2cut_369
timestamp 1717613630
transform 0 1 13427 1 0 -20073
box 16088 -7932 16222 -7868
use sky130_fd_pr__nfet_g5v0d10v5_FJGQFC  XM1 paramcells
timestamp 1717692607
transform 1 0 4664 0 1 -3159
box -357 -358 357 358
use sky130_fd_pr__pfet_g5v0d10v5_KLWMS5  XM5 paramcells
timestamp 1717691772
transform 1 0 5446 0 1 -2308
box -545 -397 545 397
use sky130_fd_pr__pfet_g5v0d10v5_KLWMS5  XM6
timestamp 1717691772
transform 1 0 6346 0 1 -2308
box -545 -397 545 397
use sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y  XM7 paramcells
timestamp 1717690002
transform 1 0 6430 0 1 -3159
box -357 -358 357 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQFS  XM8 paramcells
timestamp 1717691772
transform 1 0 5173 0 1 -3159
box -278 -358 278 358
use sky130_fd_pr__nfet_05v0_nvt_BH6ZTK  XM9 paramcells
timestamp 1717692607
transform 1 0 5762 0 1 -3159
box -437 -358 437 358
use sky130_fd_pr__nfet_g5v0d10v5_H7BQFY  XM10 paramcells
timestamp 1717691772
transform 1 0 4508 0 1 -3955
box -515 -358 515 358
use sky130_fd_pr__pfet_g5v0d10v5_AQ2WAW  XM12 paramcells
timestamp 1717690002
transform 1 0 5073 0 1 -1527
box -1809 -397 1809 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQFS  XM13
timestamp 1717691772
transform 1 0 5175 0 1 -3955
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_Z8JNCQ  XM20 paramcells
timestamp 1717691772
transform 1 0 5073 0 1 1911
box -1809 -3231 1809 3231
use sky130_fd_pr__nfet_g5v0d10v5_H7BQ24  XM22 paramcells
timestamp 1717690002
transform 1 0 6272 0 1 -3956
box -515 -358 515 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQFS  XM24
timestamp 1717691772
transform 1 0 5605 0 1 -3955
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_KLJMY6  XM25 paramcells
timestamp 1717692607
transform 1 0 3725 0 1 -2308
box -466 -397 466 397
use sky130_fd_pr__pfet_g5v0d10v5_KLWMS5  XM27
timestamp 1717691772
transform 1 0 4546 0 1 -2308
box -545 -397 545 397
use sky130_fd_pr__nfet_g5v0d10v5_UNEQFS  XM29
timestamp 1717691772
transform 1 0 4155 0 1 -3159
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_UNEQFS  XM30
timestamp 1717691772
transform 1 0 3725 0 1 -3159
box -278 -358 278 358
use sky130_fd_pr__res_xhigh_po_0p35_HLA228  XR1 paramcells
timestamp 1717716768
transform 0 1 5050 -1 0 -4833
box -367 -1748 367 1748
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XXD1 paramcells
timestamp 1717690002
transform 1 0 3634 0 1 -4088
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XXD2
timestamp 1717690002
transform 1 0 3634 0 1 -3828
box -183 -183 183 183
<< labels >>
flabel metal2 3139 4842 3339 5042 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal2 6769 -1282 6969 -1082 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal2 4034 -2396 4034 -2396 0 FreeSans 400 0 0 0 vcomp
flabel metal2 3120 -2660 3320 -2460 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal2 4884 -4077 4884 -4077 0 FreeSans 400 0 0 0 nbias
flabel metal2 3146 -3665 3346 -3465 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal2 3124 -4393 3324 -4193 0 FreeSans 256 0 0 0 ena
port 2 nsew
flabel metal1 3567 -2759 3567 -2759 0 FreeSans 400 90 0 0 pbias
flabel metal1 2863 -5640 2971 -5491 0 FreeSans 960 0 0 0 vsub
port 5 nsew
<< end >>
