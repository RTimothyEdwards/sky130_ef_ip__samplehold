magic
tech sky130A
magscale 1 2
timestamp 1717691772
<< nwell >>
rect -1809 -3231 1809 3231
<< mvpmos >>
rect -1551 2734 -1451 2934
rect -1393 2734 -1293 2934
rect -1235 2734 -1135 2934
rect -1077 2734 -977 2934
rect -919 2734 -819 2934
rect -761 2734 -661 2934
rect -603 2734 -503 2934
rect -445 2734 -345 2934
rect -287 2734 -187 2934
rect -129 2734 -29 2934
rect 29 2734 129 2934
rect 187 2734 287 2934
rect 345 2734 445 2934
rect 503 2734 603 2934
rect 661 2734 761 2934
rect 819 2734 919 2934
rect 977 2734 1077 2934
rect 1135 2734 1235 2934
rect 1293 2734 1393 2934
rect 1451 2734 1551 2934
rect -1551 2298 -1451 2498
rect -1393 2298 -1293 2498
rect -1235 2298 -1135 2498
rect -1077 2298 -977 2498
rect -919 2298 -819 2498
rect -761 2298 -661 2498
rect -603 2298 -503 2498
rect -445 2298 -345 2498
rect -287 2298 -187 2498
rect -129 2298 -29 2498
rect 29 2298 129 2498
rect 187 2298 287 2498
rect 345 2298 445 2498
rect 503 2298 603 2498
rect 661 2298 761 2498
rect 819 2298 919 2498
rect 977 2298 1077 2498
rect 1135 2298 1235 2498
rect 1293 2298 1393 2498
rect 1451 2298 1551 2498
rect -1551 1862 -1451 2062
rect -1393 1862 -1293 2062
rect -1235 1862 -1135 2062
rect -1077 1862 -977 2062
rect -919 1862 -819 2062
rect -761 1862 -661 2062
rect -603 1862 -503 2062
rect -445 1862 -345 2062
rect -287 1862 -187 2062
rect -129 1862 -29 2062
rect 29 1862 129 2062
rect 187 1862 287 2062
rect 345 1862 445 2062
rect 503 1862 603 2062
rect 661 1862 761 2062
rect 819 1862 919 2062
rect 977 1862 1077 2062
rect 1135 1862 1235 2062
rect 1293 1862 1393 2062
rect 1451 1862 1551 2062
rect -1551 1426 -1451 1626
rect -1393 1426 -1293 1626
rect -1235 1426 -1135 1626
rect -1077 1426 -977 1626
rect -919 1426 -819 1626
rect -761 1426 -661 1626
rect -603 1426 -503 1626
rect -445 1426 -345 1626
rect -287 1426 -187 1626
rect -129 1426 -29 1626
rect 29 1426 129 1626
rect 187 1426 287 1626
rect 345 1426 445 1626
rect 503 1426 603 1626
rect 661 1426 761 1626
rect 819 1426 919 1626
rect 977 1426 1077 1626
rect 1135 1426 1235 1626
rect 1293 1426 1393 1626
rect 1451 1426 1551 1626
rect -1551 990 -1451 1190
rect -1393 990 -1293 1190
rect -1235 990 -1135 1190
rect -1077 990 -977 1190
rect -919 990 -819 1190
rect -761 990 -661 1190
rect -603 990 -503 1190
rect -445 990 -345 1190
rect -287 990 -187 1190
rect -129 990 -29 1190
rect 29 990 129 1190
rect 187 990 287 1190
rect 345 990 445 1190
rect 503 990 603 1190
rect 661 990 761 1190
rect 819 990 919 1190
rect 977 990 1077 1190
rect 1135 990 1235 1190
rect 1293 990 1393 1190
rect 1451 990 1551 1190
rect -1551 554 -1451 754
rect -1393 554 -1293 754
rect -1235 554 -1135 754
rect -1077 554 -977 754
rect -919 554 -819 754
rect -761 554 -661 754
rect -603 554 -503 754
rect -445 554 -345 754
rect -287 554 -187 754
rect -129 554 -29 754
rect 29 554 129 754
rect 187 554 287 754
rect 345 554 445 754
rect 503 554 603 754
rect 661 554 761 754
rect 819 554 919 754
rect 977 554 1077 754
rect 1135 554 1235 754
rect 1293 554 1393 754
rect 1451 554 1551 754
rect -1551 118 -1451 318
rect -1393 118 -1293 318
rect -1235 118 -1135 318
rect -1077 118 -977 318
rect -919 118 -819 318
rect -761 118 -661 318
rect -603 118 -503 318
rect -445 118 -345 318
rect -287 118 -187 318
rect -129 118 -29 318
rect 29 118 129 318
rect 187 118 287 318
rect 345 118 445 318
rect 503 118 603 318
rect 661 118 761 318
rect 819 118 919 318
rect 977 118 1077 318
rect 1135 118 1235 318
rect 1293 118 1393 318
rect 1451 118 1551 318
rect -1551 -318 -1451 -118
rect -1393 -318 -1293 -118
rect -1235 -318 -1135 -118
rect -1077 -318 -977 -118
rect -919 -318 -819 -118
rect -761 -318 -661 -118
rect -603 -318 -503 -118
rect -445 -318 -345 -118
rect -287 -318 -187 -118
rect -129 -318 -29 -118
rect 29 -318 129 -118
rect 187 -318 287 -118
rect 345 -318 445 -118
rect 503 -318 603 -118
rect 661 -318 761 -118
rect 819 -318 919 -118
rect 977 -318 1077 -118
rect 1135 -318 1235 -118
rect 1293 -318 1393 -118
rect 1451 -318 1551 -118
rect -1551 -754 -1451 -554
rect -1393 -754 -1293 -554
rect -1235 -754 -1135 -554
rect -1077 -754 -977 -554
rect -919 -754 -819 -554
rect -761 -754 -661 -554
rect -603 -754 -503 -554
rect -445 -754 -345 -554
rect -287 -754 -187 -554
rect -129 -754 -29 -554
rect 29 -754 129 -554
rect 187 -754 287 -554
rect 345 -754 445 -554
rect 503 -754 603 -554
rect 661 -754 761 -554
rect 819 -754 919 -554
rect 977 -754 1077 -554
rect 1135 -754 1235 -554
rect 1293 -754 1393 -554
rect 1451 -754 1551 -554
rect -1551 -1190 -1451 -990
rect -1393 -1190 -1293 -990
rect -1235 -1190 -1135 -990
rect -1077 -1190 -977 -990
rect -919 -1190 -819 -990
rect -761 -1190 -661 -990
rect -603 -1190 -503 -990
rect -445 -1190 -345 -990
rect -287 -1190 -187 -990
rect -129 -1190 -29 -990
rect 29 -1190 129 -990
rect 187 -1190 287 -990
rect 345 -1190 445 -990
rect 503 -1190 603 -990
rect 661 -1190 761 -990
rect 819 -1190 919 -990
rect 977 -1190 1077 -990
rect 1135 -1190 1235 -990
rect 1293 -1190 1393 -990
rect 1451 -1190 1551 -990
rect -1551 -1626 -1451 -1426
rect -1393 -1626 -1293 -1426
rect -1235 -1626 -1135 -1426
rect -1077 -1626 -977 -1426
rect -919 -1626 -819 -1426
rect -761 -1626 -661 -1426
rect -603 -1626 -503 -1426
rect -445 -1626 -345 -1426
rect -287 -1626 -187 -1426
rect -129 -1626 -29 -1426
rect 29 -1626 129 -1426
rect 187 -1626 287 -1426
rect 345 -1626 445 -1426
rect 503 -1626 603 -1426
rect 661 -1626 761 -1426
rect 819 -1626 919 -1426
rect 977 -1626 1077 -1426
rect 1135 -1626 1235 -1426
rect 1293 -1626 1393 -1426
rect 1451 -1626 1551 -1426
rect -1551 -2062 -1451 -1862
rect -1393 -2062 -1293 -1862
rect -1235 -2062 -1135 -1862
rect -1077 -2062 -977 -1862
rect -919 -2062 -819 -1862
rect -761 -2062 -661 -1862
rect -603 -2062 -503 -1862
rect -445 -2062 -345 -1862
rect -287 -2062 -187 -1862
rect -129 -2062 -29 -1862
rect 29 -2062 129 -1862
rect 187 -2062 287 -1862
rect 345 -2062 445 -1862
rect 503 -2062 603 -1862
rect 661 -2062 761 -1862
rect 819 -2062 919 -1862
rect 977 -2062 1077 -1862
rect 1135 -2062 1235 -1862
rect 1293 -2062 1393 -1862
rect 1451 -2062 1551 -1862
rect -1551 -2498 -1451 -2298
rect -1393 -2498 -1293 -2298
rect -1235 -2498 -1135 -2298
rect -1077 -2498 -977 -2298
rect -919 -2498 -819 -2298
rect -761 -2498 -661 -2298
rect -603 -2498 -503 -2298
rect -445 -2498 -345 -2298
rect -287 -2498 -187 -2298
rect -129 -2498 -29 -2298
rect 29 -2498 129 -2298
rect 187 -2498 287 -2298
rect 345 -2498 445 -2298
rect 503 -2498 603 -2298
rect 661 -2498 761 -2298
rect 819 -2498 919 -2298
rect 977 -2498 1077 -2298
rect 1135 -2498 1235 -2298
rect 1293 -2498 1393 -2298
rect 1451 -2498 1551 -2298
rect -1551 -2934 -1451 -2734
rect -1393 -2934 -1293 -2734
rect -1235 -2934 -1135 -2734
rect -1077 -2934 -977 -2734
rect -919 -2934 -819 -2734
rect -761 -2934 -661 -2734
rect -603 -2934 -503 -2734
rect -445 -2934 -345 -2734
rect -287 -2934 -187 -2734
rect -129 -2934 -29 -2734
rect 29 -2934 129 -2734
rect 187 -2934 287 -2734
rect 345 -2934 445 -2734
rect 503 -2934 603 -2734
rect 661 -2934 761 -2734
rect 819 -2934 919 -2734
rect 977 -2934 1077 -2734
rect 1135 -2934 1235 -2734
rect 1293 -2934 1393 -2734
rect 1451 -2934 1551 -2734
<< mvpdiff >>
rect -1609 2922 -1551 2934
rect -1609 2746 -1597 2922
rect -1563 2746 -1551 2922
rect -1609 2734 -1551 2746
rect -1451 2922 -1393 2934
rect -1451 2746 -1439 2922
rect -1405 2746 -1393 2922
rect -1451 2734 -1393 2746
rect -1293 2922 -1235 2934
rect -1293 2746 -1281 2922
rect -1247 2746 -1235 2922
rect -1293 2734 -1235 2746
rect -1135 2922 -1077 2934
rect -1135 2746 -1123 2922
rect -1089 2746 -1077 2922
rect -1135 2734 -1077 2746
rect -977 2922 -919 2934
rect -977 2746 -965 2922
rect -931 2746 -919 2922
rect -977 2734 -919 2746
rect -819 2922 -761 2934
rect -819 2746 -807 2922
rect -773 2746 -761 2922
rect -819 2734 -761 2746
rect -661 2922 -603 2934
rect -661 2746 -649 2922
rect -615 2746 -603 2922
rect -661 2734 -603 2746
rect -503 2922 -445 2934
rect -503 2746 -491 2922
rect -457 2746 -445 2922
rect -503 2734 -445 2746
rect -345 2922 -287 2934
rect -345 2746 -333 2922
rect -299 2746 -287 2922
rect -345 2734 -287 2746
rect -187 2922 -129 2934
rect -187 2746 -175 2922
rect -141 2746 -129 2922
rect -187 2734 -129 2746
rect -29 2922 29 2934
rect -29 2746 -17 2922
rect 17 2746 29 2922
rect -29 2734 29 2746
rect 129 2922 187 2934
rect 129 2746 141 2922
rect 175 2746 187 2922
rect 129 2734 187 2746
rect 287 2922 345 2934
rect 287 2746 299 2922
rect 333 2746 345 2922
rect 287 2734 345 2746
rect 445 2922 503 2934
rect 445 2746 457 2922
rect 491 2746 503 2922
rect 445 2734 503 2746
rect 603 2922 661 2934
rect 603 2746 615 2922
rect 649 2746 661 2922
rect 603 2734 661 2746
rect 761 2922 819 2934
rect 761 2746 773 2922
rect 807 2746 819 2922
rect 761 2734 819 2746
rect 919 2922 977 2934
rect 919 2746 931 2922
rect 965 2746 977 2922
rect 919 2734 977 2746
rect 1077 2922 1135 2934
rect 1077 2746 1089 2922
rect 1123 2746 1135 2922
rect 1077 2734 1135 2746
rect 1235 2922 1293 2934
rect 1235 2746 1247 2922
rect 1281 2746 1293 2922
rect 1235 2734 1293 2746
rect 1393 2922 1451 2934
rect 1393 2746 1405 2922
rect 1439 2746 1451 2922
rect 1393 2734 1451 2746
rect 1551 2922 1609 2934
rect 1551 2746 1563 2922
rect 1597 2746 1609 2922
rect 1551 2734 1609 2746
rect -1609 2486 -1551 2498
rect -1609 2310 -1597 2486
rect -1563 2310 -1551 2486
rect -1609 2298 -1551 2310
rect -1451 2486 -1393 2498
rect -1451 2310 -1439 2486
rect -1405 2310 -1393 2486
rect -1451 2298 -1393 2310
rect -1293 2486 -1235 2498
rect -1293 2310 -1281 2486
rect -1247 2310 -1235 2486
rect -1293 2298 -1235 2310
rect -1135 2486 -1077 2498
rect -1135 2310 -1123 2486
rect -1089 2310 -1077 2486
rect -1135 2298 -1077 2310
rect -977 2486 -919 2498
rect -977 2310 -965 2486
rect -931 2310 -919 2486
rect -977 2298 -919 2310
rect -819 2486 -761 2498
rect -819 2310 -807 2486
rect -773 2310 -761 2486
rect -819 2298 -761 2310
rect -661 2486 -603 2498
rect -661 2310 -649 2486
rect -615 2310 -603 2486
rect -661 2298 -603 2310
rect -503 2486 -445 2498
rect -503 2310 -491 2486
rect -457 2310 -445 2486
rect -503 2298 -445 2310
rect -345 2486 -287 2498
rect -345 2310 -333 2486
rect -299 2310 -287 2486
rect -345 2298 -287 2310
rect -187 2486 -129 2498
rect -187 2310 -175 2486
rect -141 2310 -129 2486
rect -187 2298 -129 2310
rect -29 2486 29 2498
rect -29 2310 -17 2486
rect 17 2310 29 2486
rect -29 2298 29 2310
rect 129 2486 187 2498
rect 129 2310 141 2486
rect 175 2310 187 2486
rect 129 2298 187 2310
rect 287 2486 345 2498
rect 287 2310 299 2486
rect 333 2310 345 2486
rect 287 2298 345 2310
rect 445 2486 503 2498
rect 445 2310 457 2486
rect 491 2310 503 2486
rect 445 2298 503 2310
rect 603 2486 661 2498
rect 603 2310 615 2486
rect 649 2310 661 2486
rect 603 2298 661 2310
rect 761 2486 819 2498
rect 761 2310 773 2486
rect 807 2310 819 2486
rect 761 2298 819 2310
rect 919 2486 977 2498
rect 919 2310 931 2486
rect 965 2310 977 2486
rect 919 2298 977 2310
rect 1077 2486 1135 2498
rect 1077 2310 1089 2486
rect 1123 2310 1135 2486
rect 1077 2298 1135 2310
rect 1235 2486 1293 2498
rect 1235 2310 1247 2486
rect 1281 2310 1293 2486
rect 1235 2298 1293 2310
rect 1393 2486 1451 2498
rect 1393 2310 1405 2486
rect 1439 2310 1451 2486
rect 1393 2298 1451 2310
rect 1551 2486 1609 2498
rect 1551 2310 1563 2486
rect 1597 2310 1609 2486
rect 1551 2298 1609 2310
rect -1609 2050 -1551 2062
rect -1609 1874 -1597 2050
rect -1563 1874 -1551 2050
rect -1609 1862 -1551 1874
rect -1451 2050 -1393 2062
rect -1451 1874 -1439 2050
rect -1405 1874 -1393 2050
rect -1451 1862 -1393 1874
rect -1293 2050 -1235 2062
rect -1293 1874 -1281 2050
rect -1247 1874 -1235 2050
rect -1293 1862 -1235 1874
rect -1135 2050 -1077 2062
rect -1135 1874 -1123 2050
rect -1089 1874 -1077 2050
rect -1135 1862 -1077 1874
rect -977 2050 -919 2062
rect -977 1874 -965 2050
rect -931 1874 -919 2050
rect -977 1862 -919 1874
rect -819 2050 -761 2062
rect -819 1874 -807 2050
rect -773 1874 -761 2050
rect -819 1862 -761 1874
rect -661 2050 -603 2062
rect -661 1874 -649 2050
rect -615 1874 -603 2050
rect -661 1862 -603 1874
rect -503 2050 -445 2062
rect -503 1874 -491 2050
rect -457 1874 -445 2050
rect -503 1862 -445 1874
rect -345 2050 -287 2062
rect -345 1874 -333 2050
rect -299 1874 -287 2050
rect -345 1862 -287 1874
rect -187 2050 -129 2062
rect -187 1874 -175 2050
rect -141 1874 -129 2050
rect -187 1862 -129 1874
rect -29 2050 29 2062
rect -29 1874 -17 2050
rect 17 1874 29 2050
rect -29 1862 29 1874
rect 129 2050 187 2062
rect 129 1874 141 2050
rect 175 1874 187 2050
rect 129 1862 187 1874
rect 287 2050 345 2062
rect 287 1874 299 2050
rect 333 1874 345 2050
rect 287 1862 345 1874
rect 445 2050 503 2062
rect 445 1874 457 2050
rect 491 1874 503 2050
rect 445 1862 503 1874
rect 603 2050 661 2062
rect 603 1874 615 2050
rect 649 1874 661 2050
rect 603 1862 661 1874
rect 761 2050 819 2062
rect 761 1874 773 2050
rect 807 1874 819 2050
rect 761 1862 819 1874
rect 919 2050 977 2062
rect 919 1874 931 2050
rect 965 1874 977 2050
rect 919 1862 977 1874
rect 1077 2050 1135 2062
rect 1077 1874 1089 2050
rect 1123 1874 1135 2050
rect 1077 1862 1135 1874
rect 1235 2050 1293 2062
rect 1235 1874 1247 2050
rect 1281 1874 1293 2050
rect 1235 1862 1293 1874
rect 1393 2050 1451 2062
rect 1393 1874 1405 2050
rect 1439 1874 1451 2050
rect 1393 1862 1451 1874
rect 1551 2050 1609 2062
rect 1551 1874 1563 2050
rect 1597 1874 1609 2050
rect 1551 1862 1609 1874
rect -1609 1614 -1551 1626
rect -1609 1438 -1597 1614
rect -1563 1438 -1551 1614
rect -1609 1426 -1551 1438
rect -1451 1614 -1393 1626
rect -1451 1438 -1439 1614
rect -1405 1438 -1393 1614
rect -1451 1426 -1393 1438
rect -1293 1614 -1235 1626
rect -1293 1438 -1281 1614
rect -1247 1438 -1235 1614
rect -1293 1426 -1235 1438
rect -1135 1614 -1077 1626
rect -1135 1438 -1123 1614
rect -1089 1438 -1077 1614
rect -1135 1426 -1077 1438
rect -977 1614 -919 1626
rect -977 1438 -965 1614
rect -931 1438 -919 1614
rect -977 1426 -919 1438
rect -819 1614 -761 1626
rect -819 1438 -807 1614
rect -773 1438 -761 1614
rect -819 1426 -761 1438
rect -661 1614 -603 1626
rect -661 1438 -649 1614
rect -615 1438 -603 1614
rect -661 1426 -603 1438
rect -503 1614 -445 1626
rect -503 1438 -491 1614
rect -457 1438 -445 1614
rect -503 1426 -445 1438
rect -345 1614 -287 1626
rect -345 1438 -333 1614
rect -299 1438 -287 1614
rect -345 1426 -287 1438
rect -187 1614 -129 1626
rect -187 1438 -175 1614
rect -141 1438 -129 1614
rect -187 1426 -129 1438
rect -29 1614 29 1626
rect -29 1438 -17 1614
rect 17 1438 29 1614
rect -29 1426 29 1438
rect 129 1614 187 1626
rect 129 1438 141 1614
rect 175 1438 187 1614
rect 129 1426 187 1438
rect 287 1614 345 1626
rect 287 1438 299 1614
rect 333 1438 345 1614
rect 287 1426 345 1438
rect 445 1614 503 1626
rect 445 1438 457 1614
rect 491 1438 503 1614
rect 445 1426 503 1438
rect 603 1614 661 1626
rect 603 1438 615 1614
rect 649 1438 661 1614
rect 603 1426 661 1438
rect 761 1614 819 1626
rect 761 1438 773 1614
rect 807 1438 819 1614
rect 761 1426 819 1438
rect 919 1614 977 1626
rect 919 1438 931 1614
rect 965 1438 977 1614
rect 919 1426 977 1438
rect 1077 1614 1135 1626
rect 1077 1438 1089 1614
rect 1123 1438 1135 1614
rect 1077 1426 1135 1438
rect 1235 1614 1293 1626
rect 1235 1438 1247 1614
rect 1281 1438 1293 1614
rect 1235 1426 1293 1438
rect 1393 1614 1451 1626
rect 1393 1438 1405 1614
rect 1439 1438 1451 1614
rect 1393 1426 1451 1438
rect 1551 1614 1609 1626
rect 1551 1438 1563 1614
rect 1597 1438 1609 1614
rect 1551 1426 1609 1438
rect -1609 1178 -1551 1190
rect -1609 1002 -1597 1178
rect -1563 1002 -1551 1178
rect -1609 990 -1551 1002
rect -1451 1178 -1393 1190
rect -1451 1002 -1439 1178
rect -1405 1002 -1393 1178
rect -1451 990 -1393 1002
rect -1293 1178 -1235 1190
rect -1293 1002 -1281 1178
rect -1247 1002 -1235 1178
rect -1293 990 -1235 1002
rect -1135 1178 -1077 1190
rect -1135 1002 -1123 1178
rect -1089 1002 -1077 1178
rect -1135 990 -1077 1002
rect -977 1178 -919 1190
rect -977 1002 -965 1178
rect -931 1002 -919 1178
rect -977 990 -919 1002
rect -819 1178 -761 1190
rect -819 1002 -807 1178
rect -773 1002 -761 1178
rect -819 990 -761 1002
rect -661 1178 -603 1190
rect -661 1002 -649 1178
rect -615 1002 -603 1178
rect -661 990 -603 1002
rect -503 1178 -445 1190
rect -503 1002 -491 1178
rect -457 1002 -445 1178
rect -503 990 -445 1002
rect -345 1178 -287 1190
rect -345 1002 -333 1178
rect -299 1002 -287 1178
rect -345 990 -287 1002
rect -187 1178 -129 1190
rect -187 1002 -175 1178
rect -141 1002 -129 1178
rect -187 990 -129 1002
rect -29 1178 29 1190
rect -29 1002 -17 1178
rect 17 1002 29 1178
rect -29 990 29 1002
rect 129 1178 187 1190
rect 129 1002 141 1178
rect 175 1002 187 1178
rect 129 990 187 1002
rect 287 1178 345 1190
rect 287 1002 299 1178
rect 333 1002 345 1178
rect 287 990 345 1002
rect 445 1178 503 1190
rect 445 1002 457 1178
rect 491 1002 503 1178
rect 445 990 503 1002
rect 603 1178 661 1190
rect 603 1002 615 1178
rect 649 1002 661 1178
rect 603 990 661 1002
rect 761 1178 819 1190
rect 761 1002 773 1178
rect 807 1002 819 1178
rect 761 990 819 1002
rect 919 1178 977 1190
rect 919 1002 931 1178
rect 965 1002 977 1178
rect 919 990 977 1002
rect 1077 1178 1135 1190
rect 1077 1002 1089 1178
rect 1123 1002 1135 1178
rect 1077 990 1135 1002
rect 1235 1178 1293 1190
rect 1235 1002 1247 1178
rect 1281 1002 1293 1178
rect 1235 990 1293 1002
rect 1393 1178 1451 1190
rect 1393 1002 1405 1178
rect 1439 1002 1451 1178
rect 1393 990 1451 1002
rect 1551 1178 1609 1190
rect 1551 1002 1563 1178
rect 1597 1002 1609 1178
rect 1551 990 1609 1002
rect -1609 742 -1551 754
rect -1609 566 -1597 742
rect -1563 566 -1551 742
rect -1609 554 -1551 566
rect -1451 742 -1393 754
rect -1451 566 -1439 742
rect -1405 566 -1393 742
rect -1451 554 -1393 566
rect -1293 742 -1235 754
rect -1293 566 -1281 742
rect -1247 566 -1235 742
rect -1293 554 -1235 566
rect -1135 742 -1077 754
rect -1135 566 -1123 742
rect -1089 566 -1077 742
rect -1135 554 -1077 566
rect -977 742 -919 754
rect -977 566 -965 742
rect -931 566 -919 742
rect -977 554 -919 566
rect -819 742 -761 754
rect -819 566 -807 742
rect -773 566 -761 742
rect -819 554 -761 566
rect -661 742 -603 754
rect -661 566 -649 742
rect -615 566 -603 742
rect -661 554 -603 566
rect -503 742 -445 754
rect -503 566 -491 742
rect -457 566 -445 742
rect -503 554 -445 566
rect -345 742 -287 754
rect -345 566 -333 742
rect -299 566 -287 742
rect -345 554 -287 566
rect -187 742 -129 754
rect -187 566 -175 742
rect -141 566 -129 742
rect -187 554 -129 566
rect -29 742 29 754
rect -29 566 -17 742
rect 17 566 29 742
rect -29 554 29 566
rect 129 742 187 754
rect 129 566 141 742
rect 175 566 187 742
rect 129 554 187 566
rect 287 742 345 754
rect 287 566 299 742
rect 333 566 345 742
rect 287 554 345 566
rect 445 742 503 754
rect 445 566 457 742
rect 491 566 503 742
rect 445 554 503 566
rect 603 742 661 754
rect 603 566 615 742
rect 649 566 661 742
rect 603 554 661 566
rect 761 742 819 754
rect 761 566 773 742
rect 807 566 819 742
rect 761 554 819 566
rect 919 742 977 754
rect 919 566 931 742
rect 965 566 977 742
rect 919 554 977 566
rect 1077 742 1135 754
rect 1077 566 1089 742
rect 1123 566 1135 742
rect 1077 554 1135 566
rect 1235 742 1293 754
rect 1235 566 1247 742
rect 1281 566 1293 742
rect 1235 554 1293 566
rect 1393 742 1451 754
rect 1393 566 1405 742
rect 1439 566 1451 742
rect 1393 554 1451 566
rect 1551 742 1609 754
rect 1551 566 1563 742
rect 1597 566 1609 742
rect 1551 554 1609 566
rect -1609 306 -1551 318
rect -1609 130 -1597 306
rect -1563 130 -1551 306
rect -1609 118 -1551 130
rect -1451 306 -1393 318
rect -1451 130 -1439 306
rect -1405 130 -1393 306
rect -1451 118 -1393 130
rect -1293 306 -1235 318
rect -1293 130 -1281 306
rect -1247 130 -1235 306
rect -1293 118 -1235 130
rect -1135 306 -1077 318
rect -1135 130 -1123 306
rect -1089 130 -1077 306
rect -1135 118 -1077 130
rect -977 306 -919 318
rect -977 130 -965 306
rect -931 130 -919 306
rect -977 118 -919 130
rect -819 306 -761 318
rect -819 130 -807 306
rect -773 130 -761 306
rect -819 118 -761 130
rect -661 306 -603 318
rect -661 130 -649 306
rect -615 130 -603 306
rect -661 118 -603 130
rect -503 306 -445 318
rect -503 130 -491 306
rect -457 130 -445 306
rect -503 118 -445 130
rect -345 306 -287 318
rect -345 130 -333 306
rect -299 130 -287 306
rect -345 118 -287 130
rect -187 306 -129 318
rect -187 130 -175 306
rect -141 130 -129 306
rect -187 118 -129 130
rect -29 306 29 318
rect -29 130 -17 306
rect 17 130 29 306
rect -29 118 29 130
rect 129 306 187 318
rect 129 130 141 306
rect 175 130 187 306
rect 129 118 187 130
rect 287 306 345 318
rect 287 130 299 306
rect 333 130 345 306
rect 287 118 345 130
rect 445 306 503 318
rect 445 130 457 306
rect 491 130 503 306
rect 445 118 503 130
rect 603 306 661 318
rect 603 130 615 306
rect 649 130 661 306
rect 603 118 661 130
rect 761 306 819 318
rect 761 130 773 306
rect 807 130 819 306
rect 761 118 819 130
rect 919 306 977 318
rect 919 130 931 306
rect 965 130 977 306
rect 919 118 977 130
rect 1077 306 1135 318
rect 1077 130 1089 306
rect 1123 130 1135 306
rect 1077 118 1135 130
rect 1235 306 1293 318
rect 1235 130 1247 306
rect 1281 130 1293 306
rect 1235 118 1293 130
rect 1393 306 1451 318
rect 1393 130 1405 306
rect 1439 130 1451 306
rect 1393 118 1451 130
rect 1551 306 1609 318
rect 1551 130 1563 306
rect 1597 130 1609 306
rect 1551 118 1609 130
rect -1609 -130 -1551 -118
rect -1609 -306 -1597 -130
rect -1563 -306 -1551 -130
rect -1609 -318 -1551 -306
rect -1451 -130 -1393 -118
rect -1451 -306 -1439 -130
rect -1405 -306 -1393 -130
rect -1451 -318 -1393 -306
rect -1293 -130 -1235 -118
rect -1293 -306 -1281 -130
rect -1247 -306 -1235 -130
rect -1293 -318 -1235 -306
rect -1135 -130 -1077 -118
rect -1135 -306 -1123 -130
rect -1089 -306 -1077 -130
rect -1135 -318 -1077 -306
rect -977 -130 -919 -118
rect -977 -306 -965 -130
rect -931 -306 -919 -130
rect -977 -318 -919 -306
rect -819 -130 -761 -118
rect -819 -306 -807 -130
rect -773 -306 -761 -130
rect -819 -318 -761 -306
rect -661 -130 -603 -118
rect -661 -306 -649 -130
rect -615 -306 -603 -130
rect -661 -318 -603 -306
rect -503 -130 -445 -118
rect -503 -306 -491 -130
rect -457 -306 -445 -130
rect -503 -318 -445 -306
rect -345 -130 -287 -118
rect -345 -306 -333 -130
rect -299 -306 -287 -130
rect -345 -318 -287 -306
rect -187 -130 -129 -118
rect -187 -306 -175 -130
rect -141 -306 -129 -130
rect -187 -318 -129 -306
rect -29 -130 29 -118
rect -29 -306 -17 -130
rect 17 -306 29 -130
rect -29 -318 29 -306
rect 129 -130 187 -118
rect 129 -306 141 -130
rect 175 -306 187 -130
rect 129 -318 187 -306
rect 287 -130 345 -118
rect 287 -306 299 -130
rect 333 -306 345 -130
rect 287 -318 345 -306
rect 445 -130 503 -118
rect 445 -306 457 -130
rect 491 -306 503 -130
rect 445 -318 503 -306
rect 603 -130 661 -118
rect 603 -306 615 -130
rect 649 -306 661 -130
rect 603 -318 661 -306
rect 761 -130 819 -118
rect 761 -306 773 -130
rect 807 -306 819 -130
rect 761 -318 819 -306
rect 919 -130 977 -118
rect 919 -306 931 -130
rect 965 -306 977 -130
rect 919 -318 977 -306
rect 1077 -130 1135 -118
rect 1077 -306 1089 -130
rect 1123 -306 1135 -130
rect 1077 -318 1135 -306
rect 1235 -130 1293 -118
rect 1235 -306 1247 -130
rect 1281 -306 1293 -130
rect 1235 -318 1293 -306
rect 1393 -130 1451 -118
rect 1393 -306 1405 -130
rect 1439 -306 1451 -130
rect 1393 -318 1451 -306
rect 1551 -130 1609 -118
rect 1551 -306 1563 -130
rect 1597 -306 1609 -130
rect 1551 -318 1609 -306
rect -1609 -566 -1551 -554
rect -1609 -742 -1597 -566
rect -1563 -742 -1551 -566
rect -1609 -754 -1551 -742
rect -1451 -566 -1393 -554
rect -1451 -742 -1439 -566
rect -1405 -742 -1393 -566
rect -1451 -754 -1393 -742
rect -1293 -566 -1235 -554
rect -1293 -742 -1281 -566
rect -1247 -742 -1235 -566
rect -1293 -754 -1235 -742
rect -1135 -566 -1077 -554
rect -1135 -742 -1123 -566
rect -1089 -742 -1077 -566
rect -1135 -754 -1077 -742
rect -977 -566 -919 -554
rect -977 -742 -965 -566
rect -931 -742 -919 -566
rect -977 -754 -919 -742
rect -819 -566 -761 -554
rect -819 -742 -807 -566
rect -773 -742 -761 -566
rect -819 -754 -761 -742
rect -661 -566 -603 -554
rect -661 -742 -649 -566
rect -615 -742 -603 -566
rect -661 -754 -603 -742
rect -503 -566 -445 -554
rect -503 -742 -491 -566
rect -457 -742 -445 -566
rect -503 -754 -445 -742
rect -345 -566 -287 -554
rect -345 -742 -333 -566
rect -299 -742 -287 -566
rect -345 -754 -287 -742
rect -187 -566 -129 -554
rect -187 -742 -175 -566
rect -141 -742 -129 -566
rect -187 -754 -129 -742
rect -29 -566 29 -554
rect -29 -742 -17 -566
rect 17 -742 29 -566
rect -29 -754 29 -742
rect 129 -566 187 -554
rect 129 -742 141 -566
rect 175 -742 187 -566
rect 129 -754 187 -742
rect 287 -566 345 -554
rect 287 -742 299 -566
rect 333 -742 345 -566
rect 287 -754 345 -742
rect 445 -566 503 -554
rect 445 -742 457 -566
rect 491 -742 503 -566
rect 445 -754 503 -742
rect 603 -566 661 -554
rect 603 -742 615 -566
rect 649 -742 661 -566
rect 603 -754 661 -742
rect 761 -566 819 -554
rect 761 -742 773 -566
rect 807 -742 819 -566
rect 761 -754 819 -742
rect 919 -566 977 -554
rect 919 -742 931 -566
rect 965 -742 977 -566
rect 919 -754 977 -742
rect 1077 -566 1135 -554
rect 1077 -742 1089 -566
rect 1123 -742 1135 -566
rect 1077 -754 1135 -742
rect 1235 -566 1293 -554
rect 1235 -742 1247 -566
rect 1281 -742 1293 -566
rect 1235 -754 1293 -742
rect 1393 -566 1451 -554
rect 1393 -742 1405 -566
rect 1439 -742 1451 -566
rect 1393 -754 1451 -742
rect 1551 -566 1609 -554
rect 1551 -742 1563 -566
rect 1597 -742 1609 -566
rect 1551 -754 1609 -742
rect -1609 -1002 -1551 -990
rect -1609 -1178 -1597 -1002
rect -1563 -1178 -1551 -1002
rect -1609 -1190 -1551 -1178
rect -1451 -1002 -1393 -990
rect -1451 -1178 -1439 -1002
rect -1405 -1178 -1393 -1002
rect -1451 -1190 -1393 -1178
rect -1293 -1002 -1235 -990
rect -1293 -1178 -1281 -1002
rect -1247 -1178 -1235 -1002
rect -1293 -1190 -1235 -1178
rect -1135 -1002 -1077 -990
rect -1135 -1178 -1123 -1002
rect -1089 -1178 -1077 -1002
rect -1135 -1190 -1077 -1178
rect -977 -1002 -919 -990
rect -977 -1178 -965 -1002
rect -931 -1178 -919 -1002
rect -977 -1190 -919 -1178
rect -819 -1002 -761 -990
rect -819 -1178 -807 -1002
rect -773 -1178 -761 -1002
rect -819 -1190 -761 -1178
rect -661 -1002 -603 -990
rect -661 -1178 -649 -1002
rect -615 -1178 -603 -1002
rect -661 -1190 -603 -1178
rect -503 -1002 -445 -990
rect -503 -1178 -491 -1002
rect -457 -1178 -445 -1002
rect -503 -1190 -445 -1178
rect -345 -1002 -287 -990
rect -345 -1178 -333 -1002
rect -299 -1178 -287 -1002
rect -345 -1190 -287 -1178
rect -187 -1002 -129 -990
rect -187 -1178 -175 -1002
rect -141 -1178 -129 -1002
rect -187 -1190 -129 -1178
rect -29 -1002 29 -990
rect -29 -1178 -17 -1002
rect 17 -1178 29 -1002
rect -29 -1190 29 -1178
rect 129 -1002 187 -990
rect 129 -1178 141 -1002
rect 175 -1178 187 -1002
rect 129 -1190 187 -1178
rect 287 -1002 345 -990
rect 287 -1178 299 -1002
rect 333 -1178 345 -1002
rect 287 -1190 345 -1178
rect 445 -1002 503 -990
rect 445 -1178 457 -1002
rect 491 -1178 503 -1002
rect 445 -1190 503 -1178
rect 603 -1002 661 -990
rect 603 -1178 615 -1002
rect 649 -1178 661 -1002
rect 603 -1190 661 -1178
rect 761 -1002 819 -990
rect 761 -1178 773 -1002
rect 807 -1178 819 -1002
rect 761 -1190 819 -1178
rect 919 -1002 977 -990
rect 919 -1178 931 -1002
rect 965 -1178 977 -1002
rect 919 -1190 977 -1178
rect 1077 -1002 1135 -990
rect 1077 -1178 1089 -1002
rect 1123 -1178 1135 -1002
rect 1077 -1190 1135 -1178
rect 1235 -1002 1293 -990
rect 1235 -1178 1247 -1002
rect 1281 -1178 1293 -1002
rect 1235 -1190 1293 -1178
rect 1393 -1002 1451 -990
rect 1393 -1178 1405 -1002
rect 1439 -1178 1451 -1002
rect 1393 -1190 1451 -1178
rect 1551 -1002 1609 -990
rect 1551 -1178 1563 -1002
rect 1597 -1178 1609 -1002
rect 1551 -1190 1609 -1178
rect -1609 -1438 -1551 -1426
rect -1609 -1614 -1597 -1438
rect -1563 -1614 -1551 -1438
rect -1609 -1626 -1551 -1614
rect -1451 -1438 -1393 -1426
rect -1451 -1614 -1439 -1438
rect -1405 -1614 -1393 -1438
rect -1451 -1626 -1393 -1614
rect -1293 -1438 -1235 -1426
rect -1293 -1614 -1281 -1438
rect -1247 -1614 -1235 -1438
rect -1293 -1626 -1235 -1614
rect -1135 -1438 -1077 -1426
rect -1135 -1614 -1123 -1438
rect -1089 -1614 -1077 -1438
rect -1135 -1626 -1077 -1614
rect -977 -1438 -919 -1426
rect -977 -1614 -965 -1438
rect -931 -1614 -919 -1438
rect -977 -1626 -919 -1614
rect -819 -1438 -761 -1426
rect -819 -1614 -807 -1438
rect -773 -1614 -761 -1438
rect -819 -1626 -761 -1614
rect -661 -1438 -603 -1426
rect -661 -1614 -649 -1438
rect -615 -1614 -603 -1438
rect -661 -1626 -603 -1614
rect -503 -1438 -445 -1426
rect -503 -1614 -491 -1438
rect -457 -1614 -445 -1438
rect -503 -1626 -445 -1614
rect -345 -1438 -287 -1426
rect -345 -1614 -333 -1438
rect -299 -1614 -287 -1438
rect -345 -1626 -287 -1614
rect -187 -1438 -129 -1426
rect -187 -1614 -175 -1438
rect -141 -1614 -129 -1438
rect -187 -1626 -129 -1614
rect -29 -1438 29 -1426
rect -29 -1614 -17 -1438
rect 17 -1614 29 -1438
rect -29 -1626 29 -1614
rect 129 -1438 187 -1426
rect 129 -1614 141 -1438
rect 175 -1614 187 -1438
rect 129 -1626 187 -1614
rect 287 -1438 345 -1426
rect 287 -1614 299 -1438
rect 333 -1614 345 -1438
rect 287 -1626 345 -1614
rect 445 -1438 503 -1426
rect 445 -1614 457 -1438
rect 491 -1614 503 -1438
rect 445 -1626 503 -1614
rect 603 -1438 661 -1426
rect 603 -1614 615 -1438
rect 649 -1614 661 -1438
rect 603 -1626 661 -1614
rect 761 -1438 819 -1426
rect 761 -1614 773 -1438
rect 807 -1614 819 -1438
rect 761 -1626 819 -1614
rect 919 -1438 977 -1426
rect 919 -1614 931 -1438
rect 965 -1614 977 -1438
rect 919 -1626 977 -1614
rect 1077 -1438 1135 -1426
rect 1077 -1614 1089 -1438
rect 1123 -1614 1135 -1438
rect 1077 -1626 1135 -1614
rect 1235 -1438 1293 -1426
rect 1235 -1614 1247 -1438
rect 1281 -1614 1293 -1438
rect 1235 -1626 1293 -1614
rect 1393 -1438 1451 -1426
rect 1393 -1614 1405 -1438
rect 1439 -1614 1451 -1438
rect 1393 -1626 1451 -1614
rect 1551 -1438 1609 -1426
rect 1551 -1614 1563 -1438
rect 1597 -1614 1609 -1438
rect 1551 -1626 1609 -1614
rect -1609 -1874 -1551 -1862
rect -1609 -2050 -1597 -1874
rect -1563 -2050 -1551 -1874
rect -1609 -2062 -1551 -2050
rect -1451 -1874 -1393 -1862
rect -1451 -2050 -1439 -1874
rect -1405 -2050 -1393 -1874
rect -1451 -2062 -1393 -2050
rect -1293 -1874 -1235 -1862
rect -1293 -2050 -1281 -1874
rect -1247 -2050 -1235 -1874
rect -1293 -2062 -1235 -2050
rect -1135 -1874 -1077 -1862
rect -1135 -2050 -1123 -1874
rect -1089 -2050 -1077 -1874
rect -1135 -2062 -1077 -2050
rect -977 -1874 -919 -1862
rect -977 -2050 -965 -1874
rect -931 -2050 -919 -1874
rect -977 -2062 -919 -2050
rect -819 -1874 -761 -1862
rect -819 -2050 -807 -1874
rect -773 -2050 -761 -1874
rect -819 -2062 -761 -2050
rect -661 -1874 -603 -1862
rect -661 -2050 -649 -1874
rect -615 -2050 -603 -1874
rect -661 -2062 -603 -2050
rect -503 -1874 -445 -1862
rect -503 -2050 -491 -1874
rect -457 -2050 -445 -1874
rect -503 -2062 -445 -2050
rect -345 -1874 -287 -1862
rect -345 -2050 -333 -1874
rect -299 -2050 -287 -1874
rect -345 -2062 -287 -2050
rect -187 -1874 -129 -1862
rect -187 -2050 -175 -1874
rect -141 -2050 -129 -1874
rect -187 -2062 -129 -2050
rect -29 -1874 29 -1862
rect -29 -2050 -17 -1874
rect 17 -2050 29 -1874
rect -29 -2062 29 -2050
rect 129 -1874 187 -1862
rect 129 -2050 141 -1874
rect 175 -2050 187 -1874
rect 129 -2062 187 -2050
rect 287 -1874 345 -1862
rect 287 -2050 299 -1874
rect 333 -2050 345 -1874
rect 287 -2062 345 -2050
rect 445 -1874 503 -1862
rect 445 -2050 457 -1874
rect 491 -2050 503 -1874
rect 445 -2062 503 -2050
rect 603 -1874 661 -1862
rect 603 -2050 615 -1874
rect 649 -2050 661 -1874
rect 603 -2062 661 -2050
rect 761 -1874 819 -1862
rect 761 -2050 773 -1874
rect 807 -2050 819 -1874
rect 761 -2062 819 -2050
rect 919 -1874 977 -1862
rect 919 -2050 931 -1874
rect 965 -2050 977 -1874
rect 919 -2062 977 -2050
rect 1077 -1874 1135 -1862
rect 1077 -2050 1089 -1874
rect 1123 -2050 1135 -1874
rect 1077 -2062 1135 -2050
rect 1235 -1874 1293 -1862
rect 1235 -2050 1247 -1874
rect 1281 -2050 1293 -1874
rect 1235 -2062 1293 -2050
rect 1393 -1874 1451 -1862
rect 1393 -2050 1405 -1874
rect 1439 -2050 1451 -1874
rect 1393 -2062 1451 -2050
rect 1551 -1874 1609 -1862
rect 1551 -2050 1563 -1874
rect 1597 -2050 1609 -1874
rect 1551 -2062 1609 -2050
rect -1609 -2310 -1551 -2298
rect -1609 -2486 -1597 -2310
rect -1563 -2486 -1551 -2310
rect -1609 -2498 -1551 -2486
rect -1451 -2310 -1393 -2298
rect -1451 -2486 -1439 -2310
rect -1405 -2486 -1393 -2310
rect -1451 -2498 -1393 -2486
rect -1293 -2310 -1235 -2298
rect -1293 -2486 -1281 -2310
rect -1247 -2486 -1235 -2310
rect -1293 -2498 -1235 -2486
rect -1135 -2310 -1077 -2298
rect -1135 -2486 -1123 -2310
rect -1089 -2486 -1077 -2310
rect -1135 -2498 -1077 -2486
rect -977 -2310 -919 -2298
rect -977 -2486 -965 -2310
rect -931 -2486 -919 -2310
rect -977 -2498 -919 -2486
rect -819 -2310 -761 -2298
rect -819 -2486 -807 -2310
rect -773 -2486 -761 -2310
rect -819 -2498 -761 -2486
rect -661 -2310 -603 -2298
rect -661 -2486 -649 -2310
rect -615 -2486 -603 -2310
rect -661 -2498 -603 -2486
rect -503 -2310 -445 -2298
rect -503 -2486 -491 -2310
rect -457 -2486 -445 -2310
rect -503 -2498 -445 -2486
rect -345 -2310 -287 -2298
rect -345 -2486 -333 -2310
rect -299 -2486 -287 -2310
rect -345 -2498 -287 -2486
rect -187 -2310 -129 -2298
rect -187 -2486 -175 -2310
rect -141 -2486 -129 -2310
rect -187 -2498 -129 -2486
rect -29 -2310 29 -2298
rect -29 -2486 -17 -2310
rect 17 -2486 29 -2310
rect -29 -2498 29 -2486
rect 129 -2310 187 -2298
rect 129 -2486 141 -2310
rect 175 -2486 187 -2310
rect 129 -2498 187 -2486
rect 287 -2310 345 -2298
rect 287 -2486 299 -2310
rect 333 -2486 345 -2310
rect 287 -2498 345 -2486
rect 445 -2310 503 -2298
rect 445 -2486 457 -2310
rect 491 -2486 503 -2310
rect 445 -2498 503 -2486
rect 603 -2310 661 -2298
rect 603 -2486 615 -2310
rect 649 -2486 661 -2310
rect 603 -2498 661 -2486
rect 761 -2310 819 -2298
rect 761 -2486 773 -2310
rect 807 -2486 819 -2310
rect 761 -2498 819 -2486
rect 919 -2310 977 -2298
rect 919 -2486 931 -2310
rect 965 -2486 977 -2310
rect 919 -2498 977 -2486
rect 1077 -2310 1135 -2298
rect 1077 -2486 1089 -2310
rect 1123 -2486 1135 -2310
rect 1077 -2498 1135 -2486
rect 1235 -2310 1293 -2298
rect 1235 -2486 1247 -2310
rect 1281 -2486 1293 -2310
rect 1235 -2498 1293 -2486
rect 1393 -2310 1451 -2298
rect 1393 -2486 1405 -2310
rect 1439 -2486 1451 -2310
rect 1393 -2498 1451 -2486
rect 1551 -2310 1609 -2298
rect 1551 -2486 1563 -2310
rect 1597 -2486 1609 -2310
rect 1551 -2498 1609 -2486
rect -1609 -2746 -1551 -2734
rect -1609 -2922 -1597 -2746
rect -1563 -2922 -1551 -2746
rect -1609 -2934 -1551 -2922
rect -1451 -2746 -1393 -2734
rect -1451 -2922 -1439 -2746
rect -1405 -2922 -1393 -2746
rect -1451 -2934 -1393 -2922
rect -1293 -2746 -1235 -2734
rect -1293 -2922 -1281 -2746
rect -1247 -2922 -1235 -2746
rect -1293 -2934 -1235 -2922
rect -1135 -2746 -1077 -2734
rect -1135 -2922 -1123 -2746
rect -1089 -2922 -1077 -2746
rect -1135 -2934 -1077 -2922
rect -977 -2746 -919 -2734
rect -977 -2922 -965 -2746
rect -931 -2922 -919 -2746
rect -977 -2934 -919 -2922
rect -819 -2746 -761 -2734
rect -819 -2922 -807 -2746
rect -773 -2922 -761 -2746
rect -819 -2934 -761 -2922
rect -661 -2746 -603 -2734
rect -661 -2922 -649 -2746
rect -615 -2922 -603 -2746
rect -661 -2934 -603 -2922
rect -503 -2746 -445 -2734
rect -503 -2922 -491 -2746
rect -457 -2922 -445 -2746
rect -503 -2934 -445 -2922
rect -345 -2746 -287 -2734
rect -345 -2922 -333 -2746
rect -299 -2922 -287 -2746
rect -345 -2934 -287 -2922
rect -187 -2746 -129 -2734
rect -187 -2922 -175 -2746
rect -141 -2922 -129 -2746
rect -187 -2934 -129 -2922
rect -29 -2746 29 -2734
rect -29 -2922 -17 -2746
rect 17 -2922 29 -2746
rect -29 -2934 29 -2922
rect 129 -2746 187 -2734
rect 129 -2922 141 -2746
rect 175 -2922 187 -2746
rect 129 -2934 187 -2922
rect 287 -2746 345 -2734
rect 287 -2922 299 -2746
rect 333 -2922 345 -2746
rect 287 -2934 345 -2922
rect 445 -2746 503 -2734
rect 445 -2922 457 -2746
rect 491 -2922 503 -2746
rect 445 -2934 503 -2922
rect 603 -2746 661 -2734
rect 603 -2922 615 -2746
rect 649 -2922 661 -2746
rect 603 -2934 661 -2922
rect 761 -2746 819 -2734
rect 761 -2922 773 -2746
rect 807 -2922 819 -2746
rect 761 -2934 819 -2922
rect 919 -2746 977 -2734
rect 919 -2922 931 -2746
rect 965 -2922 977 -2746
rect 919 -2934 977 -2922
rect 1077 -2746 1135 -2734
rect 1077 -2922 1089 -2746
rect 1123 -2922 1135 -2746
rect 1077 -2934 1135 -2922
rect 1235 -2746 1293 -2734
rect 1235 -2922 1247 -2746
rect 1281 -2922 1293 -2746
rect 1235 -2934 1293 -2922
rect 1393 -2746 1451 -2734
rect 1393 -2922 1405 -2746
rect 1439 -2922 1451 -2746
rect 1393 -2934 1451 -2922
rect 1551 -2746 1609 -2734
rect 1551 -2922 1563 -2746
rect 1597 -2922 1609 -2746
rect 1551 -2934 1609 -2922
<< mvpdiffc >>
rect -1597 2746 -1563 2922
rect -1439 2746 -1405 2922
rect -1281 2746 -1247 2922
rect -1123 2746 -1089 2922
rect -965 2746 -931 2922
rect -807 2746 -773 2922
rect -649 2746 -615 2922
rect -491 2746 -457 2922
rect -333 2746 -299 2922
rect -175 2746 -141 2922
rect -17 2746 17 2922
rect 141 2746 175 2922
rect 299 2746 333 2922
rect 457 2746 491 2922
rect 615 2746 649 2922
rect 773 2746 807 2922
rect 931 2746 965 2922
rect 1089 2746 1123 2922
rect 1247 2746 1281 2922
rect 1405 2746 1439 2922
rect 1563 2746 1597 2922
rect -1597 2310 -1563 2486
rect -1439 2310 -1405 2486
rect -1281 2310 -1247 2486
rect -1123 2310 -1089 2486
rect -965 2310 -931 2486
rect -807 2310 -773 2486
rect -649 2310 -615 2486
rect -491 2310 -457 2486
rect -333 2310 -299 2486
rect -175 2310 -141 2486
rect -17 2310 17 2486
rect 141 2310 175 2486
rect 299 2310 333 2486
rect 457 2310 491 2486
rect 615 2310 649 2486
rect 773 2310 807 2486
rect 931 2310 965 2486
rect 1089 2310 1123 2486
rect 1247 2310 1281 2486
rect 1405 2310 1439 2486
rect 1563 2310 1597 2486
rect -1597 1874 -1563 2050
rect -1439 1874 -1405 2050
rect -1281 1874 -1247 2050
rect -1123 1874 -1089 2050
rect -965 1874 -931 2050
rect -807 1874 -773 2050
rect -649 1874 -615 2050
rect -491 1874 -457 2050
rect -333 1874 -299 2050
rect -175 1874 -141 2050
rect -17 1874 17 2050
rect 141 1874 175 2050
rect 299 1874 333 2050
rect 457 1874 491 2050
rect 615 1874 649 2050
rect 773 1874 807 2050
rect 931 1874 965 2050
rect 1089 1874 1123 2050
rect 1247 1874 1281 2050
rect 1405 1874 1439 2050
rect 1563 1874 1597 2050
rect -1597 1438 -1563 1614
rect -1439 1438 -1405 1614
rect -1281 1438 -1247 1614
rect -1123 1438 -1089 1614
rect -965 1438 -931 1614
rect -807 1438 -773 1614
rect -649 1438 -615 1614
rect -491 1438 -457 1614
rect -333 1438 -299 1614
rect -175 1438 -141 1614
rect -17 1438 17 1614
rect 141 1438 175 1614
rect 299 1438 333 1614
rect 457 1438 491 1614
rect 615 1438 649 1614
rect 773 1438 807 1614
rect 931 1438 965 1614
rect 1089 1438 1123 1614
rect 1247 1438 1281 1614
rect 1405 1438 1439 1614
rect 1563 1438 1597 1614
rect -1597 1002 -1563 1178
rect -1439 1002 -1405 1178
rect -1281 1002 -1247 1178
rect -1123 1002 -1089 1178
rect -965 1002 -931 1178
rect -807 1002 -773 1178
rect -649 1002 -615 1178
rect -491 1002 -457 1178
rect -333 1002 -299 1178
rect -175 1002 -141 1178
rect -17 1002 17 1178
rect 141 1002 175 1178
rect 299 1002 333 1178
rect 457 1002 491 1178
rect 615 1002 649 1178
rect 773 1002 807 1178
rect 931 1002 965 1178
rect 1089 1002 1123 1178
rect 1247 1002 1281 1178
rect 1405 1002 1439 1178
rect 1563 1002 1597 1178
rect -1597 566 -1563 742
rect -1439 566 -1405 742
rect -1281 566 -1247 742
rect -1123 566 -1089 742
rect -965 566 -931 742
rect -807 566 -773 742
rect -649 566 -615 742
rect -491 566 -457 742
rect -333 566 -299 742
rect -175 566 -141 742
rect -17 566 17 742
rect 141 566 175 742
rect 299 566 333 742
rect 457 566 491 742
rect 615 566 649 742
rect 773 566 807 742
rect 931 566 965 742
rect 1089 566 1123 742
rect 1247 566 1281 742
rect 1405 566 1439 742
rect 1563 566 1597 742
rect -1597 130 -1563 306
rect -1439 130 -1405 306
rect -1281 130 -1247 306
rect -1123 130 -1089 306
rect -965 130 -931 306
rect -807 130 -773 306
rect -649 130 -615 306
rect -491 130 -457 306
rect -333 130 -299 306
rect -175 130 -141 306
rect -17 130 17 306
rect 141 130 175 306
rect 299 130 333 306
rect 457 130 491 306
rect 615 130 649 306
rect 773 130 807 306
rect 931 130 965 306
rect 1089 130 1123 306
rect 1247 130 1281 306
rect 1405 130 1439 306
rect 1563 130 1597 306
rect -1597 -306 -1563 -130
rect -1439 -306 -1405 -130
rect -1281 -306 -1247 -130
rect -1123 -306 -1089 -130
rect -965 -306 -931 -130
rect -807 -306 -773 -130
rect -649 -306 -615 -130
rect -491 -306 -457 -130
rect -333 -306 -299 -130
rect -175 -306 -141 -130
rect -17 -306 17 -130
rect 141 -306 175 -130
rect 299 -306 333 -130
rect 457 -306 491 -130
rect 615 -306 649 -130
rect 773 -306 807 -130
rect 931 -306 965 -130
rect 1089 -306 1123 -130
rect 1247 -306 1281 -130
rect 1405 -306 1439 -130
rect 1563 -306 1597 -130
rect -1597 -742 -1563 -566
rect -1439 -742 -1405 -566
rect -1281 -742 -1247 -566
rect -1123 -742 -1089 -566
rect -965 -742 -931 -566
rect -807 -742 -773 -566
rect -649 -742 -615 -566
rect -491 -742 -457 -566
rect -333 -742 -299 -566
rect -175 -742 -141 -566
rect -17 -742 17 -566
rect 141 -742 175 -566
rect 299 -742 333 -566
rect 457 -742 491 -566
rect 615 -742 649 -566
rect 773 -742 807 -566
rect 931 -742 965 -566
rect 1089 -742 1123 -566
rect 1247 -742 1281 -566
rect 1405 -742 1439 -566
rect 1563 -742 1597 -566
rect -1597 -1178 -1563 -1002
rect -1439 -1178 -1405 -1002
rect -1281 -1178 -1247 -1002
rect -1123 -1178 -1089 -1002
rect -965 -1178 -931 -1002
rect -807 -1178 -773 -1002
rect -649 -1178 -615 -1002
rect -491 -1178 -457 -1002
rect -333 -1178 -299 -1002
rect -175 -1178 -141 -1002
rect -17 -1178 17 -1002
rect 141 -1178 175 -1002
rect 299 -1178 333 -1002
rect 457 -1178 491 -1002
rect 615 -1178 649 -1002
rect 773 -1178 807 -1002
rect 931 -1178 965 -1002
rect 1089 -1178 1123 -1002
rect 1247 -1178 1281 -1002
rect 1405 -1178 1439 -1002
rect 1563 -1178 1597 -1002
rect -1597 -1614 -1563 -1438
rect -1439 -1614 -1405 -1438
rect -1281 -1614 -1247 -1438
rect -1123 -1614 -1089 -1438
rect -965 -1614 -931 -1438
rect -807 -1614 -773 -1438
rect -649 -1614 -615 -1438
rect -491 -1614 -457 -1438
rect -333 -1614 -299 -1438
rect -175 -1614 -141 -1438
rect -17 -1614 17 -1438
rect 141 -1614 175 -1438
rect 299 -1614 333 -1438
rect 457 -1614 491 -1438
rect 615 -1614 649 -1438
rect 773 -1614 807 -1438
rect 931 -1614 965 -1438
rect 1089 -1614 1123 -1438
rect 1247 -1614 1281 -1438
rect 1405 -1614 1439 -1438
rect 1563 -1614 1597 -1438
rect -1597 -2050 -1563 -1874
rect -1439 -2050 -1405 -1874
rect -1281 -2050 -1247 -1874
rect -1123 -2050 -1089 -1874
rect -965 -2050 -931 -1874
rect -807 -2050 -773 -1874
rect -649 -2050 -615 -1874
rect -491 -2050 -457 -1874
rect -333 -2050 -299 -1874
rect -175 -2050 -141 -1874
rect -17 -2050 17 -1874
rect 141 -2050 175 -1874
rect 299 -2050 333 -1874
rect 457 -2050 491 -1874
rect 615 -2050 649 -1874
rect 773 -2050 807 -1874
rect 931 -2050 965 -1874
rect 1089 -2050 1123 -1874
rect 1247 -2050 1281 -1874
rect 1405 -2050 1439 -1874
rect 1563 -2050 1597 -1874
rect -1597 -2486 -1563 -2310
rect -1439 -2486 -1405 -2310
rect -1281 -2486 -1247 -2310
rect -1123 -2486 -1089 -2310
rect -965 -2486 -931 -2310
rect -807 -2486 -773 -2310
rect -649 -2486 -615 -2310
rect -491 -2486 -457 -2310
rect -333 -2486 -299 -2310
rect -175 -2486 -141 -2310
rect -17 -2486 17 -2310
rect 141 -2486 175 -2310
rect 299 -2486 333 -2310
rect 457 -2486 491 -2310
rect 615 -2486 649 -2310
rect 773 -2486 807 -2310
rect 931 -2486 965 -2310
rect 1089 -2486 1123 -2310
rect 1247 -2486 1281 -2310
rect 1405 -2486 1439 -2310
rect 1563 -2486 1597 -2310
rect -1597 -2922 -1563 -2746
rect -1439 -2922 -1405 -2746
rect -1281 -2922 -1247 -2746
rect -1123 -2922 -1089 -2746
rect -965 -2922 -931 -2746
rect -807 -2922 -773 -2746
rect -649 -2922 -615 -2746
rect -491 -2922 -457 -2746
rect -333 -2922 -299 -2746
rect -175 -2922 -141 -2746
rect -17 -2922 17 -2746
rect 141 -2922 175 -2746
rect 299 -2922 333 -2746
rect 457 -2922 491 -2746
rect 615 -2922 649 -2746
rect 773 -2922 807 -2746
rect 931 -2922 965 -2746
rect 1089 -2922 1123 -2746
rect 1247 -2922 1281 -2746
rect 1405 -2922 1439 -2746
rect 1563 -2922 1597 -2746
<< mvnsubdiff >>
rect -1743 3153 1743 3165
rect -1743 3119 -1635 3153
rect 1635 3119 1743 3153
rect -1743 3107 1743 3119
rect -1743 3057 -1685 3107
rect -1743 -3057 -1731 3057
rect -1697 -3057 -1685 3057
rect 1685 3057 1743 3107
rect -1743 -3107 -1685 -3057
rect 1685 -3057 1697 3057
rect 1731 -3057 1743 3057
rect 1685 -3107 1743 -3057
rect -1743 -3119 1743 -3107
rect -1743 -3153 -1635 -3119
rect 1635 -3153 1743 -3119
rect -1743 -3165 1743 -3153
<< mvnsubdiffcont >>
rect -1635 3119 1635 3153
rect -1731 -3057 -1697 3057
rect 1697 -3057 1731 3057
rect -1635 -3153 1635 -3119
<< poly >>
rect -1551 3015 -1451 3031
rect -1551 2981 -1535 3015
rect -1467 2981 -1451 3015
rect -1551 2934 -1451 2981
rect -1393 3015 -1293 3031
rect -1393 2981 -1377 3015
rect -1309 2981 -1293 3015
rect -1393 2934 -1293 2981
rect -1235 3015 -1135 3031
rect -1235 2981 -1219 3015
rect -1151 2981 -1135 3015
rect -1235 2934 -1135 2981
rect -1077 3015 -977 3031
rect -1077 2981 -1061 3015
rect -993 2981 -977 3015
rect -1077 2934 -977 2981
rect -919 3015 -819 3031
rect -919 2981 -903 3015
rect -835 2981 -819 3015
rect -919 2934 -819 2981
rect -761 3015 -661 3031
rect -761 2981 -745 3015
rect -677 2981 -661 3015
rect -761 2934 -661 2981
rect -603 3015 -503 3031
rect -603 2981 -587 3015
rect -519 2981 -503 3015
rect -603 2934 -503 2981
rect -445 3015 -345 3031
rect -445 2981 -429 3015
rect -361 2981 -345 3015
rect -445 2934 -345 2981
rect -287 3015 -187 3031
rect -287 2981 -271 3015
rect -203 2981 -187 3015
rect -287 2934 -187 2981
rect -129 3015 -29 3031
rect -129 2981 -113 3015
rect -45 2981 -29 3015
rect -129 2934 -29 2981
rect 29 3015 129 3031
rect 29 2981 45 3015
rect 113 2981 129 3015
rect 29 2934 129 2981
rect 187 3015 287 3031
rect 187 2981 203 3015
rect 271 2981 287 3015
rect 187 2934 287 2981
rect 345 3015 445 3031
rect 345 2981 361 3015
rect 429 2981 445 3015
rect 345 2934 445 2981
rect 503 3015 603 3031
rect 503 2981 519 3015
rect 587 2981 603 3015
rect 503 2934 603 2981
rect 661 3015 761 3031
rect 661 2981 677 3015
rect 745 2981 761 3015
rect 661 2934 761 2981
rect 819 3015 919 3031
rect 819 2981 835 3015
rect 903 2981 919 3015
rect 819 2934 919 2981
rect 977 3015 1077 3031
rect 977 2981 993 3015
rect 1061 2981 1077 3015
rect 977 2934 1077 2981
rect 1135 3015 1235 3031
rect 1135 2981 1151 3015
rect 1219 2981 1235 3015
rect 1135 2934 1235 2981
rect 1293 3015 1393 3031
rect 1293 2981 1309 3015
rect 1377 2981 1393 3015
rect 1293 2934 1393 2981
rect 1451 3015 1551 3031
rect 1451 2981 1467 3015
rect 1535 2981 1551 3015
rect 1451 2934 1551 2981
rect -1551 2687 -1451 2734
rect -1551 2653 -1535 2687
rect -1467 2653 -1451 2687
rect -1551 2637 -1451 2653
rect -1393 2687 -1293 2734
rect -1393 2653 -1377 2687
rect -1309 2653 -1293 2687
rect -1393 2637 -1293 2653
rect -1235 2687 -1135 2734
rect -1235 2653 -1219 2687
rect -1151 2653 -1135 2687
rect -1235 2637 -1135 2653
rect -1077 2687 -977 2734
rect -1077 2653 -1061 2687
rect -993 2653 -977 2687
rect -1077 2637 -977 2653
rect -919 2687 -819 2734
rect -919 2653 -903 2687
rect -835 2653 -819 2687
rect -919 2637 -819 2653
rect -761 2687 -661 2734
rect -761 2653 -745 2687
rect -677 2653 -661 2687
rect -761 2637 -661 2653
rect -603 2687 -503 2734
rect -603 2653 -587 2687
rect -519 2653 -503 2687
rect -603 2637 -503 2653
rect -445 2687 -345 2734
rect -445 2653 -429 2687
rect -361 2653 -345 2687
rect -445 2637 -345 2653
rect -287 2687 -187 2734
rect -287 2653 -271 2687
rect -203 2653 -187 2687
rect -287 2637 -187 2653
rect -129 2687 -29 2734
rect -129 2653 -113 2687
rect -45 2653 -29 2687
rect -129 2637 -29 2653
rect 29 2687 129 2734
rect 29 2653 45 2687
rect 113 2653 129 2687
rect 29 2637 129 2653
rect 187 2687 287 2734
rect 187 2653 203 2687
rect 271 2653 287 2687
rect 187 2637 287 2653
rect 345 2687 445 2734
rect 345 2653 361 2687
rect 429 2653 445 2687
rect 345 2637 445 2653
rect 503 2687 603 2734
rect 503 2653 519 2687
rect 587 2653 603 2687
rect 503 2637 603 2653
rect 661 2687 761 2734
rect 661 2653 677 2687
rect 745 2653 761 2687
rect 661 2637 761 2653
rect 819 2687 919 2734
rect 819 2653 835 2687
rect 903 2653 919 2687
rect 819 2637 919 2653
rect 977 2687 1077 2734
rect 977 2653 993 2687
rect 1061 2653 1077 2687
rect 977 2637 1077 2653
rect 1135 2687 1235 2734
rect 1135 2653 1151 2687
rect 1219 2653 1235 2687
rect 1135 2637 1235 2653
rect 1293 2687 1393 2734
rect 1293 2653 1309 2687
rect 1377 2653 1393 2687
rect 1293 2637 1393 2653
rect 1451 2687 1551 2734
rect 1451 2653 1467 2687
rect 1535 2653 1551 2687
rect 1451 2637 1551 2653
rect -1551 2579 -1451 2595
rect -1551 2545 -1535 2579
rect -1467 2545 -1451 2579
rect -1551 2498 -1451 2545
rect -1393 2579 -1293 2595
rect -1393 2545 -1377 2579
rect -1309 2545 -1293 2579
rect -1393 2498 -1293 2545
rect -1235 2579 -1135 2595
rect -1235 2545 -1219 2579
rect -1151 2545 -1135 2579
rect -1235 2498 -1135 2545
rect -1077 2579 -977 2595
rect -1077 2545 -1061 2579
rect -993 2545 -977 2579
rect -1077 2498 -977 2545
rect -919 2579 -819 2595
rect -919 2545 -903 2579
rect -835 2545 -819 2579
rect -919 2498 -819 2545
rect -761 2579 -661 2595
rect -761 2545 -745 2579
rect -677 2545 -661 2579
rect -761 2498 -661 2545
rect -603 2579 -503 2595
rect -603 2545 -587 2579
rect -519 2545 -503 2579
rect -603 2498 -503 2545
rect -445 2579 -345 2595
rect -445 2545 -429 2579
rect -361 2545 -345 2579
rect -445 2498 -345 2545
rect -287 2579 -187 2595
rect -287 2545 -271 2579
rect -203 2545 -187 2579
rect -287 2498 -187 2545
rect -129 2579 -29 2595
rect -129 2545 -113 2579
rect -45 2545 -29 2579
rect -129 2498 -29 2545
rect 29 2579 129 2595
rect 29 2545 45 2579
rect 113 2545 129 2579
rect 29 2498 129 2545
rect 187 2579 287 2595
rect 187 2545 203 2579
rect 271 2545 287 2579
rect 187 2498 287 2545
rect 345 2579 445 2595
rect 345 2545 361 2579
rect 429 2545 445 2579
rect 345 2498 445 2545
rect 503 2579 603 2595
rect 503 2545 519 2579
rect 587 2545 603 2579
rect 503 2498 603 2545
rect 661 2579 761 2595
rect 661 2545 677 2579
rect 745 2545 761 2579
rect 661 2498 761 2545
rect 819 2579 919 2595
rect 819 2545 835 2579
rect 903 2545 919 2579
rect 819 2498 919 2545
rect 977 2579 1077 2595
rect 977 2545 993 2579
rect 1061 2545 1077 2579
rect 977 2498 1077 2545
rect 1135 2579 1235 2595
rect 1135 2545 1151 2579
rect 1219 2545 1235 2579
rect 1135 2498 1235 2545
rect 1293 2579 1393 2595
rect 1293 2545 1309 2579
rect 1377 2545 1393 2579
rect 1293 2498 1393 2545
rect 1451 2579 1551 2595
rect 1451 2545 1467 2579
rect 1535 2545 1551 2579
rect 1451 2498 1551 2545
rect -1551 2251 -1451 2298
rect -1551 2217 -1535 2251
rect -1467 2217 -1451 2251
rect -1551 2201 -1451 2217
rect -1393 2251 -1293 2298
rect -1393 2217 -1377 2251
rect -1309 2217 -1293 2251
rect -1393 2201 -1293 2217
rect -1235 2251 -1135 2298
rect -1235 2217 -1219 2251
rect -1151 2217 -1135 2251
rect -1235 2201 -1135 2217
rect -1077 2251 -977 2298
rect -1077 2217 -1061 2251
rect -993 2217 -977 2251
rect -1077 2201 -977 2217
rect -919 2251 -819 2298
rect -919 2217 -903 2251
rect -835 2217 -819 2251
rect -919 2201 -819 2217
rect -761 2251 -661 2298
rect -761 2217 -745 2251
rect -677 2217 -661 2251
rect -761 2201 -661 2217
rect -603 2251 -503 2298
rect -603 2217 -587 2251
rect -519 2217 -503 2251
rect -603 2201 -503 2217
rect -445 2251 -345 2298
rect -445 2217 -429 2251
rect -361 2217 -345 2251
rect -445 2201 -345 2217
rect -287 2251 -187 2298
rect -287 2217 -271 2251
rect -203 2217 -187 2251
rect -287 2201 -187 2217
rect -129 2251 -29 2298
rect -129 2217 -113 2251
rect -45 2217 -29 2251
rect -129 2201 -29 2217
rect 29 2251 129 2298
rect 29 2217 45 2251
rect 113 2217 129 2251
rect 29 2201 129 2217
rect 187 2251 287 2298
rect 187 2217 203 2251
rect 271 2217 287 2251
rect 187 2201 287 2217
rect 345 2251 445 2298
rect 345 2217 361 2251
rect 429 2217 445 2251
rect 345 2201 445 2217
rect 503 2251 603 2298
rect 503 2217 519 2251
rect 587 2217 603 2251
rect 503 2201 603 2217
rect 661 2251 761 2298
rect 661 2217 677 2251
rect 745 2217 761 2251
rect 661 2201 761 2217
rect 819 2251 919 2298
rect 819 2217 835 2251
rect 903 2217 919 2251
rect 819 2201 919 2217
rect 977 2251 1077 2298
rect 977 2217 993 2251
rect 1061 2217 1077 2251
rect 977 2201 1077 2217
rect 1135 2251 1235 2298
rect 1135 2217 1151 2251
rect 1219 2217 1235 2251
rect 1135 2201 1235 2217
rect 1293 2251 1393 2298
rect 1293 2217 1309 2251
rect 1377 2217 1393 2251
rect 1293 2201 1393 2217
rect 1451 2251 1551 2298
rect 1451 2217 1467 2251
rect 1535 2217 1551 2251
rect 1451 2201 1551 2217
rect -1551 2143 -1451 2159
rect -1551 2109 -1535 2143
rect -1467 2109 -1451 2143
rect -1551 2062 -1451 2109
rect -1393 2143 -1293 2159
rect -1393 2109 -1377 2143
rect -1309 2109 -1293 2143
rect -1393 2062 -1293 2109
rect -1235 2143 -1135 2159
rect -1235 2109 -1219 2143
rect -1151 2109 -1135 2143
rect -1235 2062 -1135 2109
rect -1077 2143 -977 2159
rect -1077 2109 -1061 2143
rect -993 2109 -977 2143
rect -1077 2062 -977 2109
rect -919 2143 -819 2159
rect -919 2109 -903 2143
rect -835 2109 -819 2143
rect -919 2062 -819 2109
rect -761 2143 -661 2159
rect -761 2109 -745 2143
rect -677 2109 -661 2143
rect -761 2062 -661 2109
rect -603 2143 -503 2159
rect -603 2109 -587 2143
rect -519 2109 -503 2143
rect -603 2062 -503 2109
rect -445 2143 -345 2159
rect -445 2109 -429 2143
rect -361 2109 -345 2143
rect -445 2062 -345 2109
rect -287 2143 -187 2159
rect -287 2109 -271 2143
rect -203 2109 -187 2143
rect -287 2062 -187 2109
rect -129 2143 -29 2159
rect -129 2109 -113 2143
rect -45 2109 -29 2143
rect -129 2062 -29 2109
rect 29 2143 129 2159
rect 29 2109 45 2143
rect 113 2109 129 2143
rect 29 2062 129 2109
rect 187 2143 287 2159
rect 187 2109 203 2143
rect 271 2109 287 2143
rect 187 2062 287 2109
rect 345 2143 445 2159
rect 345 2109 361 2143
rect 429 2109 445 2143
rect 345 2062 445 2109
rect 503 2143 603 2159
rect 503 2109 519 2143
rect 587 2109 603 2143
rect 503 2062 603 2109
rect 661 2143 761 2159
rect 661 2109 677 2143
rect 745 2109 761 2143
rect 661 2062 761 2109
rect 819 2143 919 2159
rect 819 2109 835 2143
rect 903 2109 919 2143
rect 819 2062 919 2109
rect 977 2143 1077 2159
rect 977 2109 993 2143
rect 1061 2109 1077 2143
rect 977 2062 1077 2109
rect 1135 2143 1235 2159
rect 1135 2109 1151 2143
rect 1219 2109 1235 2143
rect 1135 2062 1235 2109
rect 1293 2143 1393 2159
rect 1293 2109 1309 2143
rect 1377 2109 1393 2143
rect 1293 2062 1393 2109
rect 1451 2143 1551 2159
rect 1451 2109 1467 2143
rect 1535 2109 1551 2143
rect 1451 2062 1551 2109
rect -1551 1815 -1451 1862
rect -1551 1781 -1535 1815
rect -1467 1781 -1451 1815
rect -1551 1765 -1451 1781
rect -1393 1815 -1293 1862
rect -1393 1781 -1377 1815
rect -1309 1781 -1293 1815
rect -1393 1765 -1293 1781
rect -1235 1815 -1135 1862
rect -1235 1781 -1219 1815
rect -1151 1781 -1135 1815
rect -1235 1765 -1135 1781
rect -1077 1815 -977 1862
rect -1077 1781 -1061 1815
rect -993 1781 -977 1815
rect -1077 1765 -977 1781
rect -919 1815 -819 1862
rect -919 1781 -903 1815
rect -835 1781 -819 1815
rect -919 1765 -819 1781
rect -761 1815 -661 1862
rect -761 1781 -745 1815
rect -677 1781 -661 1815
rect -761 1765 -661 1781
rect -603 1815 -503 1862
rect -603 1781 -587 1815
rect -519 1781 -503 1815
rect -603 1765 -503 1781
rect -445 1815 -345 1862
rect -445 1781 -429 1815
rect -361 1781 -345 1815
rect -445 1765 -345 1781
rect -287 1815 -187 1862
rect -287 1781 -271 1815
rect -203 1781 -187 1815
rect -287 1765 -187 1781
rect -129 1815 -29 1862
rect -129 1781 -113 1815
rect -45 1781 -29 1815
rect -129 1765 -29 1781
rect 29 1815 129 1862
rect 29 1781 45 1815
rect 113 1781 129 1815
rect 29 1765 129 1781
rect 187 1815 287 1862
rect 187 1781 203 1815
rect 271 1781 287 1815
rect 187 1765 287 1781
rect 345 1815 445 1862
rect 345 1781 361 1815
rect 429 1781 445 1815
rect 345 1765 445 1781
rect 503 1815 603 1862
rect 503 1781 519 1815
rect 587 1781 603 1815
rect 503 1765 603 1781
rect 661 1815 761 1862
rect 661 1781 677 1815
rect 745 1781 761 1815
rect 661 1765 761 1781
rect 819 1815 919 1862
rect 819 1781 835 1815
rect 903 1781 919 1815
rect 819 1765 919 1781
rect 977 1815 1077 1862
rect 977 1781 993 1815
rect 1061 1781 1077 1815
rect 977 1765 1077 1781
rect 1135 1815 1235 1862
rect 1135 1781 1151 1815
rect 1219 1781 1235 1815
rect 1135 1765 1235 1781
rect 1293 1815 1393 1862
rect 1293 1781 1309 1815
rect 1377 1781 1393 1815
rect 1293 1765 1393 1781
rect 1451 1815 1551 1862
rect 1451 1781 1467 1815
rect 1535 1781 1551 1815
rect 1451 1765 1551 1781
rect -1551 1707 -1451 1723
rect -1551 1673 -1535 1707
rect -1467 1673 -1451 1707
rect -1551 1626 -1451 1673
rect -1393 1707 -1293 1723
rect -1393 1673 -1377 1707
rect -1309 1673 -1293 1707
rect -1393 1626 -1293 1673
rect -1235 1707 -1135 1723
rect -1235 1673 -1219 1707
rect -1151 1673 -1135 1707
rect -1235 1626 -1135 1673
rect -1077 1707 -977 1723
rect -1077 1673 -1061 1707
rect -993 1673 -977 1707
rect -1077 1626 -977 1673
rect -919 1707 -819 1723
rect -919 1673 -903 1707
rect -835 1673 -819 1707
rect -919 1626 -819 1673
rect -761 1707 -661 1723
rect -761 1673 -745 1707
rect -677 1673 -661 1707
rect -761 1626 -661 1673
rect -603 1707 -503 1723
rect -603 1673 -587 1707
rect -519 1673 -503 1707
rect -603 1626 -503 1673
rect -445 1707 -345 1723
rect -445 1673 -429 1707
rect -361 1673 -345 1707
rect -445 1626 -345 1673
rect -287 1707 -187 1723
rect -287 1673 -271 1707
rect -203 1673 -187 1707
rect -287 1626 -187 1673
rect -129 1707 -29 1723
rect -129 1673 -113 1707
rect -45 1673 -29 1707
rect -129 1626 -29 1673
rect 29 1707 129 1723
rect 29 1673 45 1707
rect 113 1673 129 1707
rect 29 1626 129 1673
rect 187 1707 287 1723
rect 187 1673 203 1707
rect 271 1673 287 1707
rect 187 1626 287 1673
rect 345 1707 445 1723
rect 345 1673 361 1707
rect 429 1673 445 1707
rect 345 1626 445 1673
rect 503 1707 603 1723
rect 503 1673 519 1707
rect 587 1673 603 1707
rect 503 1626 603 1673
rect 661 1707 761 1723
rect 661 1673 677 1707
rect 745 1673 761 1707
rect 661 1626 761 1673
rect 819 1707 919 1723
rect 819 1673 835 1707
rect 903 1673 919 1707
rect 819 1626 919 1673
rect 977 1707 1077 1723
rect 977 1673 993 1707
rect 1061 1673 1077 1707
rect 977 1626 1077 1673
rect 1135 1707 1235 1723
rect 1135 1673 1151 1707
rect 1219 1673 1235 1707
rect 1135 1626 1235 1673
rect 1293 1707 1393 1723
rect 1293 1673 1309 1707
rect 1377 1673 1393 1707
rect 1293 1626 1393 1673
rect 1451 1707 1551 1723
rect 1451 1673 1467 1707
rect 1535 1673 1551 1707
rect 1451 1626 1551 1673
rect -1551 1379 -1451 1426
rect -1551 1345 -1535 1379
rect -1467 1345 -1451 1379
rect -1551 1329 -1451 1345
rect -1393 1379 -1293 1426
rect -1393 1345 -1377 1379
rect -1309 1345 -1293 1379
rect -1393 1329 -1293 1345
rect -1235 1379 -1135 1426
rect -1235 1345 -1219 1379
rect -1151 1345 -1135 1379
rect -1235 1329 -1135 1345
rect -1077 1379 -977 1426
rect -1077 1345 -1061 1379
rect -993 1345 -977 1379
rect -1077 1329 -977 1345
rect -919 1379 -819 1426
rect -919 1345 -903 1379
rect -835 1345 -819 1379
rect -919 1329 -819 1345
rect -761 1379 -661 1426
rect -761 1345 -745 1379
rect -677 1345 -661 1379
rect -761 1329 -661 1345
rect -603 1379 -503 1426
rect -603 1345 -587 1379
rect -519 1345 -503 1379
rect -603 1329 -503 1345
rect -445 1379 -345 1426
rect -445 1345 -429 1379
rect -361 1345 -345 1379
rect -445 1329 -345 1345
rect -287 1379 -187 1426
rect -287 1345 -271 1379
rect -203 1345 -187 1379
rect -287 1329 -187 1345
rect -129 1379 -29 1426
rect -129 1345 -113 1379
rect -45 1345 -29 1379
rect -129 1329 -29 1345
rect 29 1379 129 1426
rect 29 1345 45 1379
rect 113 1345 129 1379
rect 29 1329 129 1345
rect 187 1379 287 1426
rect 187 1345 203 1379
rect 271 1345 287 1379
rect 187 1329 287 1345
rect 345 1379 445 1426
rect 345 1345 361 1379
rect 429 1345 445 1379
rect 345 1329 445 1345
rect 503 1379 603 1426
rect 503 1345 519 1379
rect 587 1345 603 1379
rect 503 1329 603 1345
rect 661 1379 761 1426
rect 661 1345 677 1379
rect 745 1345 761 1379
rect 661 1329 761 1345
rect 819 1379 919 1426
rect 819 1345 835 1379
rect 903 1345 919 1379
rect 819 1329 919 1345
rect 977 1379 1077 1426
rect 977 1345 993 1379
rect 1061 1345 1077 1379
rect 977 1329 1077 1345
rect 1135 1379 1235 1426
rect 1135 1345 1151 1379
rect 1219 1345 1235 1379
rect 1135 1329 1235 1345
rect 1293 1379 1393 1426
rect 1293 1345 1309 1379
rect 1377 1345 1393 1379
rect 1293 1329 1393 1345
rect 1451 1379 1551 1426
rect 1451 1345 1467 1379
rect 1535 1345 1551 1379
rect 1451 1329 1551 1345
rect -1551 1271 -1451 1287
rect -1551 1237 -1535 1271
rect -1467 1237 -1451 1271
rect -1551 1190 -1451 1237
rect -1393 1271 -1293 1287
rect -1393 1237 -1377 1271
rect -1309 1237 -1293 1271
rect -1393 1190 -1293 1237
rect -1235 1271 -1135 1287
rect -1235 1237 -1219 1271
rect -1151 1237 -1135 1271
rect -1235 1190 -1135 1237
rect -1077 1271 -977 1287
rect -1077 1237 -1061 1271
rect -993 1237 -977 1271
rect -1077 1190 -977 1237
rect -919 1271 -819 1287
rect -919 1237 -903 1271
rect -835 1237 -819 1271
rect -919 1190 -819 1237
rect -761 1271 -661 1287
rect -761 1237 -745 1271
rect -677 1237 -661 1271
rect -761 1190 -661 1237
rect -603 1271 -503 1287
rect -603 1237 -587 1271
rect -519 1237 -503 1271
rect -603 1190 -503 1237
rect -445 1271 -345 1287
rect -445 1237 -429 1271
rect -361 1237 -345 1271
rect -445 1190 -345 1237
rect -287 1271 -187 1287
rect -287 1237 -271 1271
rect -203 1237 -187 1271
rect -287 1190 -187 1237
rect -129 1271 -29 1287
rect -129 1237 -113 1271
rect -45 1237 -29 1271
rect -129 1190 -29 1237
rect 29 1271 129 1287
rect 29 1237 45 1271
rect 113 1237 129 1271
rect 29 1190 129 1237
rect 187 1271 287 1287
rect 187 1237 203 1271
rect 271 1237 287 1271
rect 187 1190 287 1237
rect 345 1271 445 1287
rect 345 1237 361 1271
rect 429 1237 445 1271
rect 345 1190 445 1237
rect 503 1271 603 1287
rect 503 1237 519 1271
rect 587 1237 603 1271
rect 503 1190 603 1237
rect 661 1271 761 1287
rect 661 1237 677 1271
rect 745 1237 761 1271
rect 661 1190 761 1237
rect 819 1271 919 1287
rect 819 1237 835 1271
rect 903 1237 919 1271
rect 819 1190 919 1237
rect 977 1271 1077 1287
rect 977 1237 993 1271
rect 1061 1237 1077 1271
rect 977 1190 1077 1237
rect 1135 1271 1235 1287
rect 1135 1237 1151 1271
rect 1219 1237 1235 1271
rect 1135 1190 1235 1237
rect 1293 1271 1393 1287
rect 1293 1237 1309 1271
rect 1377 1237 1393 1271
rect 1293 1190 1393 1237
rect 1451 1271 1551 1287
rect 1451 1237 1467 1271
rect 1535 1237 1551 1271
rect 1451 1190 1551 1237
rect -1551 943 -1451 990
rect -1551 909 -1535 943
rect -1467 909 -1451 943
rect -1551 893 -1451 909
rect -1393 943 -1293 990
rect -1393 909 -1377 943
rect -1309 909 -1293 943
rect -1393 893 -1293 909
rect -1235 943 -1135 990
rect -1235 909 -1219 943
rect -1151 909 -1135 943
rect -1235 893 -1135 909
rect -1077 943 -977 990
rect -1077 909 -1061 943
rect -993 909 -977 943
rect -1077 893 -977 909
rect -919 943 -819 990
rect -919 909 -903 943
rect -835 909 -819 943
rect -919 893 -819 909
rect -761 943 -661 990
rect -761 909 -745 943
rect -677 909 -661 943
rect -761 893 -661 909
rect -603 943 -503 990
rect -603 909 -587 943
rect -519 909 -503 943
rect -603 893 -503 909
rect -445 943 -345 990
rect -445 909 -429 943
rect -361 909 -345 943
rect -445 893 -345 909
rect -287 943 -187 990
rect -287 909 -271 943
rect -203 909 -187 943
rect -287 893 -187 909
rect -129 943 -29 990
rect -129 909 -113 943
rect -45 909 -29 943
rect -129 893 -29 909
rect 29 943 129 990
rect 29 909 45 943
rect 113 909 129 943
rect 29 893 129 909
rect 187 943 287 990
rect 187 909 203 943
rect 271 909 287 943
rect 187 893 287 909
rect 345 943 445 990
rect 345 909 361 943
rect 429 909 445 943
rect 345 893 445 909
rect 503 943 603 990
rect 503 909 519 943
rect 587 909 603 943
rect 503 893 603 909
rect 661 943 761 990
rect 661 909 677 943
rect 745 909 761 943
rect 661 893 761 909
rect 819 943 919 990
rect 819 909 835 943
rect 903 909 919 943
rect 819 893 919 909
rect 977 943 1077 990
rect 977 909 993 943
rect 1061 909 1077 943
rect 977 893 1077 909
rect 1135 943 1235 990
rect 1135 909 1151 943
rect 1219 909 1235 943
rect 1135 893 1235 909
rect 1293 943 1393 990
rect 1293 909 1309 943
rect 1377 909 1393 943
rect 1293 893 1393 909
rect 1451 943 1551 990
rect 1451 909 1467 943
rect 1535 909 1551 943
rect 1451 893 1551 909
rect -1551 835 -1451 851
rect -1551 801 -1535 835
rect -1467 801 -1451 835
rect -1551 754 -1451 801
rect -1393 835 -1293 851
rect -1393 801 -1377 835
rect -1309 801 -1293 835
rect -1393 754 -1293 801
rect -1235 835 -1135 851
rect -1235 801 -1219 835
rect -1151 801 -1135 835
rect -1235 754 -1135 801
rect -1077 835 -977 851
rect -1077 801 -1061 835
rect -993 801 -977 835
rect -1077 754 -977 801
rect -919 835 -819 851
rect -919 801 -903 835
rect -835 801 -819 835
rect -919 754 -819 801
rect -761 835 -661 851
rect -761 801 -745 835
rect -677 801 -661 835
rect -761 754 -661 801
rect -603 835 -503 851
rect -603 801 -587 835
rect -519 801 -503 835
rect -603 754 -503 801
rect -445 835 -345 851
rect -445 801 -429 835
rect -361 801 -345 835
rect -445 754 -345 801
rect -287 835 -187 851
rect -287 801 -271 835
rect -203 801 -187 835
rect -287 754 -187 801
rect -129 835 -29 851
rect -129 801 -113 835
rect -45 801 -29 835
rect -129 754 -29 801
rect 29 835 129 851
rect 29 801 45 835
rect 113 801 129 835
rect 29 754 129 801
rect 187 835 287 851
rect 187 801 203 835
rect 271 801 287 835
rect 187 754 287 801
rect 345 835 445 851
rect 345 801 361 835
rect 429 801 445 835
rect 345 754 445 801
rect 503 835 603 851
rect 503 801 519 835
rect 587 801 603 835
rect 503 754 603 801
rect 661 835 761 851
rect 661 801 677 835
rect 745 801 761 835
rect 661 754 761 801
rect 819 835 919 851
rect 819 801 835 835
rect 903 801 919 835
rect 819 754 919 801
rect 977 835 1077 851
rect 977 801 993 835
rect 1061 801 1077 835
rect 977 754 1077 801
rect 1135 835 1235 851
rect 1135 801 1151 835
rect 1219 801 1235 835
rect 1135 754 1235 801
rect 1293 835 1393 851
rect 1293 801 1309 835
rect 1377 801 1393 835
rect 1293 754 1393 801
rect 1451 835 1551 851
rect 1451 801 1467 835
rect 1535 801 1551 835
rect 1451 754 1551 801
rect -1551 507 -1451 554
rect -1551 473 -1535 507
rect -1467 473 -1451 507
rect -1551 457 -1451 473
rect -1393 507 -1293 554
rect -1393 473 -1377 507
rect -1309 473 -1293 507
rect -1393 457 -1293 473
rect -1235 507 -1135 554
rect -1235 473 -1219 507
rect -1151 473 -1135 507
rect -1235 457 -1135 473
rect -1077 507 -977 554
rect -1077 473 -1061 507
rect -993 473 -977 507
rect -1077 457 -977 473
rect -919 507 -819 554
rect -919 473 -903 507
rect -835 473 -819 507
rect -919 457 -819 473
rect -761 507 -661 554
rect -761 473 -745 507
rect -677 473 -661 507
rect -761 457 -661 473
rect -603 507 -503 554
rect -603 473 -587 507
rect -519 473 -503 507
rect -603 457 -503 473
rect -445 507 -345 554
rect -445 473 -429 507
rect -361 473 -345 507
rect -445 457 -345 473
rect -287 507 -187 554
rect -287 473 -271 507
rect -203 473 -187 507
rect -287 457 -187 473
rect -129 507 -29 554
rect -129 473 -113 507
rect -45 473 -29 507
rect -129 457 -29 473
rect 29 507 129 554
rect 29 473 45 507
rect 113 473 129 507
rect 29 457 129 473
rect 187 507 287 554
rect 187 473 203 507
rect 271 473 287 507
rect 187 457 287 473
rect 345 507 445 554
rect 345 473 361 507
rect 429 473 445 507
rect 345 457 445 473
rect 503 507 603 554
rect 503 473 519 507
rect 587 473 603 507
rect 503 457 603 473
rect 661 507 761 554
rect 661 473 677 507
rect 745 473 761 507
rect 661 457 761 473
rect 819 507 919 554
rect 819 473 835 507
rect 903 473 919 507
rect 819 457 919 473
rect 977 507 1077 554
rect 977 473 993 507
rect 1061 473 1077 507
rect 977 457 1077 473
rect 1135 507 1235 554
rect 1135 473 1151 507
rect 1219 473 1235 507
rect 1135 457 1235 473
rect 1293 507 1393 554
rect 1293 473 1309 507
rect 1377 473 1393 507
rect 1293 457 1393 473
rect 1451 507 1551 554
rect 1451 473 1467 507
rect 1535 473 1551 507
rect 1451 457 1551 473
rect -1551 399 -1451 415
rect -1551 365 -1535 399
rect -1467 365 -1451 399
rect -1551 318 -1451 365
rect -1393 399 -1293 415
rect -1393 365 -1377 399
rect -1309 365 -1293 399
rect -1393 318 -1293 365
rect -1235 399 -1135 415
rect -1235 365 -1219 399
rect -1151 365 -1135 399
rect -1235 318 -1135 365
rect -1077 399 -977 415
rect -1077 365 -1061 399
rect -993 365 -977 399
rect -1077 318 -977 365
rect -919 399 -819 415
rect -919 365 -903 399
rect -835 365 -819 399
rect -919 318 -819 365
rect -761 399 -661 415
rect -761 365 -745 399
rect -677 365 -661 399
rect -761 318 -661 365
rect -603 399 -503 415
rect -603 365 -587 399
rect -519 365 -503 399
rect -603 318 -503 365
rect -445 399 -345 415
rect -445 365 -429 399
rect -361 365 -345 399
rect -445 318 -345 365
rect -287 399 -187 415
rect -287 365 -271 399
rect -203 365 -187 399
rect -287 318 -187 365
rect -129 399 -29 415
rect -129 365 -113 399
rect -45 365 -29 399
rect -129 318 -29 365
rect 29 399 129 415
rect 29 365 45 399
rect 113 365 129 399
rect 29 318 129 365
rect 187 399 287 415
rect 187 365 203 399
rect 271 365 287 399
rect 187 318 287 365
rect 345 399 445 415
rect 345 365 361 399
rect 429 365 445 399
rect 345 318 445 365
rect 503 399 603 415
rect 503 365 519 399
rect 587 365 603 399
rect 503 318 603 365
rect 661 399 761 415
rect 661 365 677 399
rect 745 365 761 399
rect 661 318 761 365
rect 819 399 919 415
rect 819 365 835 399
rect 903 365 919 399
rect 819 318 919 365
rect 977 399 1077 415
rect 977 365 993 399
rect 1061 365 1077 399
rect 977 318 1077 365
rect 1135 399 1235 415
rect 1135 365 1151 399
rect 1219 365 1235 399
rect 1135 318 1235 365
rect 1293 399 1393 415
rect 1293 365 1309 399
rect 1377 365 1393 399
rect 1293 318 1393 365
rect 1451 399 1551 415
rect 1451 365 1467 399
rect 1535 365 1551 399
rect 1451 318 1551 365
rect -1551 71 -1451 118
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1551 21 -1451 37
rect -1393 71 -1293 118
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1393 21 -1293 37
rect -1235 71 -1135 118
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1235 21 -1135 37
rect -1077 71 -977 118
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -1077 21 -977 37
rect -919 71 -819 118
rect -919 37 -903 71
rect -835 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 118
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 118
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 118
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 118
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 118
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 118
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 118
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 118
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect 819 71 919 118
rect 819 37 835 71
rect 903 37 919 71
rect 819 21 919 37
rect 977 71 1077 118
rect 977 37 993 71
rect 1061 37 1077 71
rect 977 21 1077 37
rect 1135 71 1235 118
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1135 21 1235 37
rect 1293 71 1393 118
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1293 21 1393 37
rect 1451 71 1551 118
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1451 21 1551 37
rect -1551 -37 -1451 -21
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1551 -118 -1451 -71
rect -1393 -37 -1293 -21
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1393 -118 -1293 -71
rect -1235 -37 -1135 -21
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1235 -118 -1135 -71
rect -1077 -37 -977 -21
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -1077 -118 -977 -71
rect -919 -37 -819 -21
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -919 -118 -819 -71
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -118 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -118 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -118 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -118 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -118 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -118 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -118 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -118 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -118 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -118 761 -71
rect 819 -37 919 -21
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 819 -118 919 -71
rect 977 -37 1077 -21
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 977 -118 1077 -71
rect 1135 -37 1235 -21
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1135 -118 1235 -71
rect 1293 -37 1393 -21
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1293 -118 1393 -71
rect 1451 -37 1551 -21
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1451 -118 1551 -71
rect -1551 -365 -1451 -318
rect -1551 -399 -1535 -365
rect -1467 -399 -1451 -365
rect -1551 -415 -1451 -399
rect -1393 -365 -1293 -318
rect -1393 -399 -1377 -365
rect -1309 -399 -1293 -365
rect -1393 -415 -1293 -399
rect -1235 -365 -1135 -318
rect -1235 -399 -1219 -365
rect -1151 -399 -1135 -365
rect -1235 -415 -1135 -399
rect -1077 -365 -977 -318
rect -1077 -399 -1061 -365
rect -993 -399 -977 -365
rect -1077 -415 -977 -399
rect -919 -365 -819 -318
rect -919 -399 -903 -365
rect -835 -399 -819 -365
rect -919 -415 -819 -399
rect -761 -365 -661 -318
rect -761 -399 -745 -365
rect -677 -399 -661 -365
rect -761 -415 -661 -399
rect -603 -365 -503 -318
rect -603 -399 -587 -365
rect -519 -399 -503 -365
rect -603 -415 -503 -399
rect -445 -365 -345 -318
rect -445 -399 -429 -365
rect -361 -399 -345 -365
rect -445 -415 -345 -399
rect -287 -365 -187 -318
rect -287 -399 -271 -365
rect -203 -399 -187 -365
rect -287 -415 -187 -399
rect -129 -365 -29 -318
rect -129 -399 -113 -365
rect -45 -399 -29 -365
rect -129 -415 -29 -399
rect 29 -365 129 -318
rect 29 -399 45 -365
rect 113 -399 129 -365
rect 29 -415 129 -399
rect 187 -365 287 -318
rect 187 -399 203 -365
rect 271 -399 287 -365
rect 187 -415 287 -399
rect 345 -365 445 -318
rect 345 -399 361 -365
rect 429 -399 445 -365
rect 345 -415 445 -399
rect 503 -365 603 -318
rect 503 -399 519 -365
rect 587 -399 603 -365
rect 503 -415 603 -399
rect 661 -365 761 -318
rect 661 -399 677 -365
rect 745 -399 761 -365
rect 661 -415 761 -399
rect 819 -365 919 -318
rect 819 -399 835 -365
rect 903 -399 919 -365
rect 819 -415 919 -399
rect 977 -365 1077 -318
rect 977 -399 993 -365
rect 1061 -399 1077 -365
rect 977 -415 1077 -399
rect 1135 -365 1235 -318
rect 1135 -399 1151 -365
rect 1219 -399 1235 -365
rect 1135 -415 1235 -399
rect 1293 -365 1393 -318
rect 1293 -399 1309 -365
rect 1377 -399 1393 -365
rect 1293 -415 1393 -399
rect 1451 -365 1551 -318
rect 1451 -399 1467 -365
rect 1535 -399 1551 -365
rect 1451 -415 1551 -399
rect -1551 -473 -1451 -457
rect -1551 -507 -1535 -473
rect -1467 -507 -1451 -473
rect -1551 -554 -1451 -507
rect -1393 -473 -1293 -457
rect -1393 -507 -1377 -473
rect -1309 -507 -1293 -473
rect -1393 -554 -1293 -507
rect -1235 -473 -1135 -457
rect -1235 -507 -1219 -473
rect -1151 -507 -1135 -473
rect -1235 -554 -1135 -507
rect -1077 -473 -977 -457
rect -1077 -507 -1061 -473
rect -993 -507 -977 -473
rect -1077 -554 -977 -507
rect -919 -473 -819 -457
rect -919 -507 -903 -473
rect -835 -507 -819 -473
rect -919 -554 -819 -507
rect -761 -473 -661 -457
rect -761 -507 -745 -473
rect -677 -507 -661 -473
rect -761 -554 -661 -507
rect -603 -473 -503 -457
rect -603 -507 -587 -473
rect -519 -507 -503 -473
rect -603 -554 -503 -507
rect -445 -473 -345 -457
rect -445 -507 -429 -473
rect -361 -507 -345 -473
rect -445 -554 -345 -507
rect -287 -473 -187 -457
rect -287 -507 -271 -473
rect -203 -507 -187 -473
rect -287 -554 -187 -507
rect -129 -473 -29 -457
rect -129 -507 -113 -473
rect -45 -507 -29 -473
rect -129 -554 -29 -507
rect 29 -473 129 -457
rect 29 -507 45 -473
rect 113 -507 129 -473
rect 29 -554 129 -507
rect 187 -473 287 -457
rect 187 -507 203 -473
rect 271 -507 287 -473
rect 187 -554 287 -507
rect 345 -473 445 -457
rect 345 -507 361 -473
rect 429 -507 445 -473
rect 345 -554 445 -507
rect 503 -473 603 -457
rect 503 -507 519 -473
rect 587 -507 603 -473
rect 503 -554 603 -507
rect 661 -473 761 -457
rect 661 -507 677 -473
rect 745 -507 761 -473
rect 661 -554 761 -507
rect 819 -473 919 -457
rect 819 -507 835 -473
rect 903 -507 919 -473
rect 819 -554 919 -507
rect 977 -473 1077 -457
rect 977 -507 993 -473
rect 1061 -507 1077 -473
rect 977 -554 1077 -507
rect 1135 -473 1235 -457
rect 1135 -507 1151 -473
rect 1219 -507 1235 -473
rect 1135 -554 1235 -507
rect 1293 -473 1393 -457
rect 1293 -507 1309 -473
rect 1377 -507 1393 -473
rect 1293 -554 1393 -507
rect 1451 -473 1551 -457
rect 1451 -507 1467 -473
rect 1535 -507 1551 -473
rect 1451 -554 1551 -507
rect -1551 -801 -1451 -754
rect -1551 -835 -1535 -801
rect -1467 -835 -1451 -801
rect -1551 -851 -1451 -835
rect -1393 -801 -1293 -754
rect -1393 -835 -1377 -801
rect -1309 -835 -1293 -801
rect -1393 -851 -1293 -835
rect -1235 -801 -1135 -754
rect -1235 -835 -1219 -801
rect -1151 -835 -1135 -801
rect -1235 -851 -1135 -835
rect -1077 -801 -977 -754
rect -1077 -835 -1061 -801
rect -993 -835 -977 -801
rect -1077 -851 -977 -835
rect -919 -801 -819 -754
rect -919 -835 -903 -801
rect -835 -835 -819 -801
rect -919 -851 -819 -835
rect -761 -801 -661 -754
rect -761 -835 -745 -801
rect -677 -835 -661 -801
rect -761 -851 -661 -835
rect -603 -801 -503 -754
rect -603 -835 -587 -801
rect -519 -835 -503 -801
rect -603 -851 -503 -835
rect -445 -801 -345 -754
rect -445 -835 -429 -801
rect -361 -835 -345 -801
rect -445 -851 -345 -835
rect -287 -801 -187 -754
rect -287 -835 -271 -801
rect -203 -835 -187 -801
rect -287 -851 -187 -835
rect -129 -801 -29 -754
rect -129 -835 -113 -801
rect -45 -835 -29 -801
rect -129 -851 -29 -835
rect 29 -801 129 -754
rect 29 -835 45 -801
rect 113 -835 129 -801
rect 29 -851 129 -835
rect 187 -801 287 -754
rect 187 -835 203 -801
rect 271 -835 287 -801
rect 187 -851 287 -835
rect 345 -801 445 -754
rect 345 -835 361 -801
rect 429 -835 445 -801
rect 345 -851 445 -835
rect 503 -801 603 -754
rect 503 -835 519 -801
rect 587 -835 603 -801
rect 503 -851 603 -835
rect 661 -801 761 -754
rect 661 -835 677 -801
rect 745 -835 761 -801
rect 661 -851 761 -835
rect 819 -801 919 -754
rect 819 -835 835 -801
rect 903 -835 919 -801
rect 819 -851 919 -835
rect 977 -801 1077 -754
rect 977 -835 993 -801
rect 1061 -835 1077 -801
rect 977 -851 1077 -835
rect 1135 -801 1235 -754
rect 1135 -835 1151 -801
rect 1219 -835 1235 -801
rect 1135 -851 1235 -835
rect 1293 -801 1393 -754
rect 1293 -835 1309 -801
rect 1377 -835 1393 -801
rect 1293 -851 1393 -835
rect 1451 -801 1551 -754
rect 1451 -835 1467 -801
rect 1535 -835 1551 -801
rect 1451 -851 1551 -835
rect -1551 -909 -1451 -893
rect -1551 -943 -1535 -909
rect -1467 -943 -1451 -909
rect -1551 -990 -1451 -943
rect -1393 -909 -1293 -893
rect -1393 -943 -1377 -909
rect -1309 -943 -1293 -909
rect -1393 -990 -1293 -943
rect -1235 -909 -1135 -893
rect -1235 -943 -1219 -909
rect -1151 -943 -1135 -909
rect -1235 -990 -1135 -943
rect -1077 -909 -977 -893
rect -1077 -943 -1061 -909
rect -993 -943 -977 -909
rect -1077 -990 -977 -943
rect -919 -909 -819 -893
rect -919 -943 -903 -909
rect -835 -943 -819 -909
rect -919 -990 -819 -943
rect -761 -909 -661 -893
rect -761 -943 -745 -909
rect -677 -943 -661 -909
rect -761 -990 -661 -943
rect -603 -909 -503 -893
rect -603 -943 -587 -909
rect -519 -943 -503 -909
rect -603 -990 -503 -943
rect -445 -909 -345 -893
rect -445 -943 -429 -909
rect -361 -943 -345 -909
rect -445 -990 -345 -943
rect -287 -909 -187 -893
rect -287 -943 -271 -909
rect -203 -943 -187 -909
rect -287 -990 -187 -943
rect -129 -909 -29 -893
rect -129 -943 -113 -909
rect -45 -943 -29 -909
rect -129 -990 -29 -943
rect 29 -909 129 -893
rect 29 -943 45 -909
rect 113 -943 129 -909
rect 29 -990 129 -943
rect 187 -909 287 -893
rect 187 -943 203 -909
rect 271 -943 287 -909
rect 187 -990 287 -943
rect 345 -909 445 -893
rect 345 -943 361 -909
rect 429 -943 445 -909
rect 345 -990 445 -943
rect 503 -909 603 -893
rect 503 -943 519 -909
rect 587 -943 603 -909
rect 503 -990 603 -943
rect 661 -909 761 -893
rect 661 -943 677 -909
rect 745 -943 761 -909
rect 661 -990 761 -943
rect 819 -909 919 -893
rect 819 -943 835 -909
rect 903 -943 919 -909
rect 819 -990 919 -943
rect 977 -909 1077 -893
rect 977 -943 993 -909
rect 1061 -943 1077 -909
rect 977 -990 1077 -943
rect 1135 -909 1235 -893
rect 1135 -943 1151 -909
rect 1219 -943 1235 -909
rect 1135 -990 1235 -943
rect 1293 -909 1393 -893
rect 1293 -943 1309 -909
rect 1377 -943 1393 -909
rect 1293 -990 1393 -943
rect 1451 -909 1551 -893
rect 1451 -943 1467 -909
rect 1535 -943 1551 -909
rect 1451 -990 1551 -943
rect -1551 -1237 -1451 -1190
rect -1551 -1271 -1535 -1237
rect -1467 -1271 -1451 -1237
rect -1551 -1287 -1451 -1271
rect -1393 -1237 -1293 -1190
rect -1393 -1271 -1377 -1237
rect -1309 -1271 -1293 -1237
rect -1393 -1287 -1293 -1271
rect -1235 -1237 -1135 -1190
rect -1235 -1271 -1219 -1237
rect -1151 -1271 -1135 -1237
rect -1235 -1287 -1135 -1271
rect -1077 -1237 -977 -1190
rect -1077 -1271 -1061 -1237
rect -993 -1271 -977 -1237
rect -1077 -1287 -977 -1271
rect -919 -1237 -819 -1190
rect -919 -1271 -903 -1237
rect -835 -1271 -819 -1237
rect -919 -1287 -819 -1271
rect -761 -1237 -661 -1190
rect -761 -1271 -745 -1237
rect -677 -1271 -661 -1237
rect -761 -1287 -661 -1271
rect -603 -1237 -503 -1190
rect -603 -1271 -587 -1237
rect -519 -1271 -503 -1237
rect -603 -1287 -503 -1271
rect -445 -1237 -345 -1190
rect -445 -1271 -429 -1237
rect -361 -1271 -345 -1237
rect -445 -1287 -345 -1271
rect -287 -1237 -187 -1190
rect -287 -1271 -271 -1237
rect -203 -1271 -187 -1237
rect -287 -1287 -187 -1271
rect -129 -1237 -29 -1190
rect -129 -1271 -113 -1237
rect -45 -1271 -29 -1237
rect -129 -1287 -29 -1271
rect 29 -1237 129 -1190
rect 29 -1271 45 -1237
rect 113 -1271 129 -1237
rect 29 -1287 129 -1271
rect 187 -1237 287 -1190
rect 187 -1271 203 -1237
rect 271 -1271 287 -1237
rect 187 -1287 287 -1271
rect 345 -1237 445 -1190
rect 345 -1271 361 -1237
rect 429 -1271 445 -1237
rect 345 -1287 445 -1271
rect 503 -1237 603 -1190
rect 503 -1271 519 -1237
rect 587 -1271 603 -1237
rect 503 -1287 603 -1271
rect 661 -1237 761 -1190
rect 661 -1271 677 -1237
rect 745 -1271 761 -1237
rect 661 -1287 761 -1271
rect 819 -1237 919 -1190
rect 819 -1271 835 -1237
rect 903 -1271 919 -1237
rect 819 -1287 919 -1271
rect 977 -1237 1077 -1190
rect 977 -1271 993 -1237
rect 1061 -1271 1077 -1237
rect 977 -1287 1077 -1271
rect 1135 -1237 1235 -1190
rect 1135 -1271 1151 -1237
rect 1219 -1271 1235 -1237
rect 1135 -1287 1235 -1271
rect 1293 -1237 1393 -1190
rect 1293 -1271 1309 -1237
rect 1377 -1271 1393 -1237
rect 1293 -1287 1393 -1271
rect 1451 -1237 1551 -1190
rect 1451 -1271 1467 -1237
rect 1535 -1271 1551 -1237
rect 1451 -1287 1551 -1271
rect -1551 -1345 -1451 -1329
rect -1551 -1379 -1535 -1345
rect -1467 -1379 -1451 -1345
rect -1551 -1426 -1451 -1379
rect -1393 -1345 -1293 -1329
rect -1393 -1379 -1377 -1345
rect -1309 -1379 -1293 -1345
rect -1393 -1426 -1293 -1379
rect -1235 -1345 -1135 -1329
rect -1235 -1379 -1219 -1345
rect -1151 -1379 -1135 -1345
rect -1235 -1426 -1135 -1379
rect -1077 -1345 -977 -1329
rect -1077 -1379 -1061 -1345
rect -993 -1379 -977 -1345
rect -1077 -1426 -977 -1379
rect -919 -1345 -819 -1329
rect -919 -1379 -903 -1345
rect -835 -1379 -819 -1345
rect -919 -1426 -819 -1379
rect -761 -1345 -661 -1329
rect -761 -1379 -745 -1345
rect -677 -1379 -661 -1345
rect -761 -1426 -661 -1379
rect -603 -1345 -503 -1329
rect -603 -1379 -587 -1345
rect -519 -1379 -503 -1345
rect -603 -1426 -503 -1379
rect -445 -1345 -345 -1329
rect -445 -1379 -429 -1345
rect -361 -1379 -345 -1345
rect -445 -1426 -345 -1379
rect -287 -1345 -187 -1329
rect -287 -1379 -271 -1345
rect -203 -1379 -187 -1345
rect -287 -1426 -187 -1379
rect -129 -1345 -29 -1329
rect -129 -1379 -113 -1345
rect -45 -1379 -29 -1345
rect -129 -1426 -29 -1379
rect 29 -1345 129 -1329
rect 29 -1379 45 -1345
rect 113 -1379 129 -1345
rect 29 -1426 129 -1379
rect 187 -1345 287 -1329
rect 187 -1379 203 -1345
rect 271 -1379 287 -1345
rect 187 -1426 287 -1379
rect 345 -1345 445 -1329
rect 345 -1379 361 -1345
rect 429 -1379 445 -1345
rect 345 -1426 445 -1379
rect 503 -1345 603 -1329
rect 503 -1379 519 -1345
rect 587 -1379 603 -1345
rect 503 -1426 603 -1379
rect 661 -1345 761 -1329
rect 661 -1379 677 -1345
rect 745 -1379 761 -1345
rect 661 -1426 761 -1379
rect 819 -1345 919 -1329
rect 819 -1379 835 -1345
rect 903 -1379 919 -1345
rect 819 -1426 919 -1379
rect 977 -1345 1077 -1329
rect 977 -1379 993 -1345
rect 1061 -1379 1077 -1345
rect 977 -1426 1077 -1379
rect 1135 -1345 1235 -1329
rect 1135 -1379 1151 -1345
rect 1219 -1379 1235 -1345
rect 1135 -1426 1235 -1379
rect 1293 -1345 1393 -1329
rect 1293 -1379 1309 -1345
rect 1377 -1379 1393 -1345
rect 1293 -1426 1393 -1379
rect 1451 -1345 1551 -1329
rect 1451 -1379 1467 -1345
rect 1535 -1379 1551 -1345
rect 1451 -1426 1551 -1379
rect -1551 -1673 -1451 -1626
rect -1551 -1707 -1535 -1673
rect -1467 -1707 -1451 -1673
rect -1551 -1723 -1451 -1707
rect -1393 -1673 -1293 -1626
rect -1393 -1707 -1377 -1673
rect -1309 -1707 -1293 -1673
rect -1393 -1723 -1293 -1707
rect -1235 -1673 -1135 -1626
rect -1235 -1707 -1219 -1673
rect -1151 -1707 -1135 -1673
rect -1235 -1723 -1135 -1707
rect -1077 -1673 -977 -1626
rect -1077 -1707 -1061 -1673
rect -993 -1707 -977 -1673
rect -1077 -1723 -977 -1707
rect -919 -1673 -819 -1626
rect -919 -1707 -903 -1673
rect -835 -1707 -819 -1673
rect -919 -1723 -819 -1707
rect -761 -1673 -661 -1626
rect -761 -1707 -745 -1673
rect -677 -1707 -661 -1673
rect -761 -1723 -661 -1707
rect -603 -1673 -503 -1626
rect -603 -1707 -587 -1673
rect -519 -1707 -503 -1673
rect -603 -1723 -503 -1707
rect -445 -1673 -345 -1626
rect -445 -1707 -429 -1673
rect -361 -1707 -345 -1673
rect -445 -1723 -345 -1707
rect -287 -1673 -187 -1626
rect -287 -1707 -271 -1673
rect -203 -1707 -187 -1673
rect -287 -1723 -187 -1707
rect -129 -1673 -29 -1626
rect -129 -1707 -113 -1673
rect -45 -1707 -29 -1673
rect -129 -1723 -29 -1707
rect 29 -1673 129 -1626
rect 29 -1707 45 -1673
rect 113 -1707 129 -1673
rect 29 -1723 129 -1707
rect 187 -1673 287 -1626
rect 187 -1707 203 -1673
rect 271 -1707 287 -1673
rect 187 -1723 287 -1707
rect 345 -1673 445 -1626
rect 345 -1707 361 -1673
rect 429 -1707 445 -1673
rect 345 -1723 445 -1707
rect 503 -1673 603 -1626
rect 503 -1707 519 -1673
rect 587 -1707 603 -1673
rect 503 -1723 603 -1707
rect 661 -1673 761 -1626
rect 661 -1707 677 -1673
rect 745 -1707 761 -1673
rect 661 -1723 761 -1707
rect 819 -1673 919 -1626
rect 819 -1707 835 -1673
rect 903 -1707 919 -1673
rect 819 -1723 919 -1707
rect 977 -1673 1077 -1626
rect 977 -1707 993 -1673
rect 1061 -1707 1077 -1673
rect 977 -1723 1077 -1707
rect 1135 -1673 1235 -1626
rect 1135 -1707 1151 -1673
rect 1219 -1707 1235 -1673
rect 1135 -1723 1235 -1707
rect 1293 -1673 1393 -1626
rect 1293 -1707 1309 -1673
rect 1377 -1707 1393 -1673
rect 1293 -1723 1393 -1707
rect 1451 -1673 1551 -1626
rect 1451 -1707 1467 -1673
rect 1535 -1707 1551 -1673
rect 1451 -1723 1551 -1707
rect -1551 -1781 -1451 -1765
rect -1551 -1815 -1535 -1781
rect -1467 -1815 -1451 -1781
rect -1551 -1862 -1451 -1815
rect -1393 -1781 -1293 -1765
rect -1393 -1815 -1377 -1781
rect -1309 -1815 -1293 -1781
rect -1393 -1862 -1293 -1815
rect -1235 -1781 -1135 -1765
rect -1235 -1815 -1219 -1781
rect -1151 -1815 -1135 -1781
rect -1235 -1862 -1135 -1815
rect -1077 -1781 -977 -1765
rect -1077 -1815 -1061 -1781
rect -993 -1815 -977 -1781
rect -1077 -1862 -977 -1815
rect -919 -1781 -819 -1765
rect -919 -1815 -903 -1781
rect -835 -1815 -819 -1781
rect -919 -1862 -819 -1815
rect -761 -1781 -661 -1765
rect -761 -1815 -745 -1781
rect -677 -1815 -661 -1781
rect -761 -1862 -661 -1815
rect -603 -1781 -503 -1765
rect -603 -1815 -587 -1781
rect -519 -1815 -503 -1781
rect -603 -1862 -503 -1815
rect -445 -1781 -345 -1765
rect -445 -1815 -429 -1781
rect -361 -1815 -345 -1781
rect -445 -1862 -345 -1815
rect -287 -1781 -187 -1765
rect -287 -1815 -271 -1781
rect -203 -1815 -187 -1781
rect -287 -1862 -187 -1815
rect -129 -1781 -29 -1765
rect -129 -1815 -113 -1781
rect -45 -1815 -29 -1781
rect -129 -1862 -29 -1815
rect 29 -1781 129 -1765
rect 29 -1815 45 -1781
rect 113 -1815 129 -1781
rect 29 -1862 129 -1815
rect 187 -1781 287 -1765
rect 187 -1815 203 -1781
rect 271 -1815 287 -1781
rect 187 -1862 287 -1815
rect 345 -1781 445 -1765
rect 345 -1815 361 -1781
rect 429 -1815 445 -1781
rect 345 -1862 445 -1815
rect 503 -1781 603 -1765
rect 503 -1815 519 -1781
rect 587 -1815 603 -1781
rect 503 -1862 603 -1815
rect 661 -1781 761 -1765
rect 661 -1815 677 -1781
rect 745 -1815 761 -1781
rect 661 -1862 761 -1815
rect 819 -1781 919 -1765
rect 819 -1815 835 -1781
rect 903 -1815 919 -1781
rect 819 -1862 919 -1815
rect 977 -1781 1077 -1765
rect 977 -1815 993 -1781
rect 1061 -1815 1077 -1781
rect 977 -1862 1077 -1815
rect 1135 -1781 1235 -1765
rect 1135 -1815 1151 -1781
rect 1219 -1815 1235 -1781
rect 1135 -1862 1235 -1815
rect 1293 -1781 1393 -1765
rect 1293 -1815 1309 -1781
rect 1377 -1815 1393 -1781
rect 1293 -1862 1393 -1815
rect 1451 -1781 1551 -1765
rect 1451 -1815 1467 -1781
rect 1535 -1815 1551 -1781
rect 1451 -1862 1551 -1815
rect -1551 -2109 -1451 -2062
rect -1551 -2143 -1535 -2109
rect -1467 -2143 -1451 -2109
rect -1551 -2159 -1451 -2143
rect -1393 -2109 -1293 -2062
rect -1393 -2143 -1377 -2109
rect -1309 -2143 -1293 -2109
rect -1393 -2159 -1293 -2143
rect -1235 -2109 -1135 -2062
rect -1235 -2143 -1219 -2109
rect -1151 -2143 -1135 -2109
rect -1235 -2159 -1135 -2143
rect -1077 -2109 -977 -2062
rect -1077 -2143 -1061 -2109
rect -993 -2143 -977 -2109
rect -1077 -2159 -977 -2143
rect -919 -2109 -819 -2062
rect -919 -2143 -903 -2109
rect -835 -2143 -819 -2109
rect -919 -2159 -819 -2143
rect -761 -2109 -661 -2062
rect -761 -2143 -745 -2109
rect -677 -2143 -661 -2109
rect -761 -2159 -661 -2143
rect -603 -2109 -503 -2062
rect -603 -2143 -587 -2109
rect -519 -2143 -503 -2109
rect -603 -2159 -503 -2143
rect -445 -2109 -345 -2062
rect -445 -2143 -429 -2109
rect -361 -2143 -345 -2109
rect -445 -2159 -345 -2143
rect -287 -2109 -187 -2062
rect -287 -2143 -271 -2109
rect -203 -2143 -187 -2109
rect -287 -2159 -187 -2143
rect -129 -2109 -29 -2062
rect -129 -2143 -113 -2109
rect -45 -2143 -29 -2109
rect -129 -2159 -29 -2143
rect 29 -2109 129 -2062
rect 29 -2143 45 -2109
rect 113 -2143 129 -2109
rect 29 -2159 129 -2143
rect 187 -2109 287 -2062
rect 187 -2143 203 -2109
rect 271 -2143 287 -2109
rect 187 -2159 287 -2143
rect 345 -2109 445 -2062
rect 345 -2143 361 -2109
rect 429 -2143 445 -2109
rect 345 -2159 445 -2143
rect 503 -2109 603 -2062
rect 503 -2143 519 -2109
rect 587 -2143 603 -2109
rect 503 -2159 603 -2143
rect 661 -2109 761 -2062
rect 661 -2143 677 -2109
rect 745 -2143 761 -2109
rect 661 -2159 761 -2143
rect 819 -2109 919 -2062
rect 819 -2143 835 -2109
rect 903 -2143 919 -2109
rect 819 -2159 919 -2143
rect 977 -2109 1077 -2062
rect 977 -2143 993 -2109
rect 1061 -2143 1077 -2109
rect 977 -2159 1077 -2143
rect 1135 -2109 1235 -2062
rect 1135 -2143 1151 -2109
rect 1219 -2143 1235 -2109
rect 1135 -2159 1235 -2143
rect 1293 -2109 1393 -2062
rect 1293 -2143 1309 -2109
rect 1377 -2143 1393 -2109
rect 1293 -2159 1393 -2143
rect 1451 -2109 1551 -2062
rect 1451 -2143 1467 -2109
rect 1535 -2143 1551 -2109
rect 1451 -2159 1551 -2143
rect -1551 -2217 -1451 -2201
rect -1551 -2251 -1535 -2217
rect -1467 -2251 -1451 -2217
rect -1551 -2298 -1451 -2251
rect -1393 -2217 -1293 -2201
rect -1393 -2251 -1377 -2217
rect -1309 -2251 -1293 -2217
rect -1393 -2298 -1293 -2251
rect -1235 -2217 -1135 -2201
rect -1235 -2251 -1219 -2217
rect -1151 -2251 -1135 -2217
rect -1235 -2298 -1135 -2251
rect -1077 -2217 -977 -2201
rect -1077 -2251 -1061 -2217
rect -993 -2251 -977 -2217
rect -1077 -2298 -977 -2251
rect -919 -2217 -819 -2201
rect -919 -2251 -903 -2217
rect -835 -2251 -819 -2217
rect -919 -2298 -819 -2251
rect -761 -2217 -661 -2201
rect -761 -2251 -745 -2217
rect -677 -2251 -661 -2217
rect -761 -2298 -661 -2251
rect -603 -2217 -503 -2201
rect -603 -2251 -587 -2217
rect -519 -2251 -503 -2217
rect -603 -2298 -503 -2251
rect -445 -2217 -345 -2201
rect -445 -2251 -429 -2217
rect -361 -2251 -345 -2217
rect -445 -2298 -345 -2251
rect -287 -2217 -187 -2201
rect -287 -2251 -271 -2217
rect -203 -2251 -187 -2217
rect -287 -2298 -187 -2251
rect -129 -2217 -29 -2201
rect -129 -2251 -113 -2217
rect -45 -2251 -29 -2217
rect -129 -2298 -29 -2251
rect 29 -2217 129 -2201
rect 29 -2251 45 -2217
rect 113 -2251 129 -2217
rect 29 -2298 129 -2251
rect 187 -2217 287 -2201
rect 187 -2251 203 -2217
rect 271 -2251 287 -2217
rect 187 -2298 287 -2251
rect 345 -2217 445 -2201
rect 345 -2251 361 -2217
rect 429 -2251 445 -2217
rect 345 -2298 445 -2251
rect 503 -2217 603 -2201
rect 503 -2251 519 -2217
rect 587 -2251 603 -2217
rect 503 -2298 603 -2251
rect 661 -2217 761 -2201
rect 661 -2251 677 -2217
rect 745 -2251 761 -2217
rect 661 -2298 761 -2251
rect 819 -2217 919 -2201
rect 819 -2251 835 -2217
rect 903 -2251 919 -2217
rect 819 -2298 919 -2251
rect 977 -2217 1077 -2201
rect 977 -2251 993 -2217
rect 1061 -2251 1077 -2217
rect 977 -2298 1077 -2251
rect 1135 -2217 1235 -2201
rect 1135 -2251 1151 -2217
rect 1219 -2251 1235 -2217
rect 1135 -2298 1235 -2251
rect 1293 -2217 1393 -2201
rect 1293 -2251 1309 -2217
rect 1377 -2251 1393 -2217
rect 1293 -2298 1393 -2251
rect 1451 -2217 1551 -2201
rect 1451 -2251 1467 -2217
rect 1535 -2251 1551 -2217
rect 1451 -2298 1551 -2251
rect -1551 -2545 -1451 -2498
rect -1551 -2579 -1535 -2545
rect -1467 -2579 -1451 -2545
rect -1551 -2595 -1451 -2579
rect -1393 -2545 -1293 -2498
rect -1393 -2579 -1377 -2545
rect -1309 -2579 -1293 -2545
rect -1393 -2595 -1293 -2579
rect -1235 -2545 -1135 -2498
rect -1235 -2579 -1219 -2545
rect -1151 -2579 -1135 -2545
rect -1235 -2595 -1135 -2579
rect -1077 -2545 -977 -2498
rect -1077 -2579 -1061 -2545
rect -993 -2579 -977 -2545
rect -1077 -2595 -977 -2579
rect -919 -2545 -819 -2498
rect -919 -2579 -903 -2545
rect -835 -2579 -819 -2545
rect -919 -2595 -819 -2579
rect -761 -2545 -661 -2498
rect -761 -2579 -745 -2545
rect -677 -2579 -661 -2545
rect -761 -2595 -661 -2579
rect -603 -2545 -503 -2498
rect -603 -2579 -587 -2545
rect -519 -2579 -503 -2545
rect -603 -2595 -503 -2579
rect -445 -2545 -345 -2498
rect -445 -2579 -429 -2545
rect -361 -2579 -345 -2545
rect -445 -2595 -345 -2579
rect -287 -2545 -187 -2498
rect -287 -2579 -271 -2545
rect -203 -2579 -187 -2545
rect -287 -2595 -187 -2579
rect -129 -2545 -29 -2498
rect -129 -2579 -113 -2545
rect -45 -2579 -29 -2545
rect -129 -2595 -29 -2579
rect 29 -2545 129 -2498
rect 29 -2579 45 -2545
rect 113 -2579 129 -2545
rect 29 -2595 129 -2579
rect 187 -2545 287 -2498
rect 187 -2579 203 -2545
rect 271 -2579 287 -2545
rect 187 -2595 287 -2579
rect 345 -2545 445 -2498
rect 345 -2579 361 -2545
rect 429 -2579 445 -2545
rect 345 -2595 445 -2579
rect 503 -2545 603 -2498
rect 503 -2579 519 -2545
rect 587 -2579 603 -2545
rect 503 -2595 603 -2579
rect 661 -2545 761 -2498
rect 661 -2579 677 -2545
rect 745 -2579 761 -2545
rect 661 -2595 761 -2579
rect 819 -2545 919 -2498
rect 819 -2579 835 -2545
rect 903 -2579 919 -2545
rect 819 -2595 919 -2579
rect 977 -2545 1077 -2498
rect 977 -2579 993 -2545
rect 1061 -2579 1077 -2545
rect 977 -2595 1077 -2579
rect 1135 -2545 1235 -2498
rect 1135 -2579 1151 -2545
rect 1219 -2579 1235 -2545
rect 1135 -2595 1235 -2579
rect 1293 -2545 1393 -2498
rect 1293 -2579 1309 -2545
rect 1377 -2579 1393 -2545
rect 1293 -2595 1393 -2579
rect 1451 -2545 1551 -2498
rect 1451 -2579 1467 -2545
rect 1535 -2579 1551 -2545
rect 1451 -2595 1551 -2579
rect -1551 -2653 -1451 -2637
rect -1551 -2687 -1535 -2653
rect -1467 -2687 -1451 -2653
rect -1551 -2734 -1451 -2687
rect -1393 -2653 -1293 -2637
rect -1393 -2687 -1377 -2653
rect -1309 -2687 -1293 -2653
rect -1393 -2734 -1293 -2687
rect -1235 -2653 -1135 -2637
rect -1235 -2687 -1219 -2653
rect -1151 -2687 -1135 -2653
rect -1235 -2734 -1135 -2687
rect -1077 -2653 -977 -2637
rect -1077 -2687 -1061 -2653
rect -993 -2687 -977 -2653
rect -1077 -2734 -977 -2687
rect -919 -2653 -819 -2637
rect -919 -2687 -903 -2653
rect -835 -2687 -819 -2653
rect -919 -2734 -819 -2687
rect -761 -2653 -661 -2637
rect -761 -2687 -745 -2653
rect -677 -2687 -661 -2653
rect -761 -2734 -661 -2687
rect -603 -2653 -503 -2637
rect -603 -2687 -587 -2653
rect -519 -2687 -503 -2653
rect -603 -2734 -503 -2687
rect -445 -2653 -345 -2637
rect -445 -2687 -429 -2653
rect -361 -2687 -345 -2653
rect -445 -2734 -345 -2687
rect -287 -2653 -187 -2637
rect -287 -2687 -271 -2653
rect -203 -2687 -187 -2653
rect -287 -2734 -187 -2687
rect -129 -2653 -29 -2637
rect -129 -2687 -113 -2653
rect -45 -2687 -29 -2653
rect -129 -2734 -29 -2687
rect 29 -2653 129 -2637
rect 29 -2687 45 -2653
rect 113 -2687 129 -2653
rect 29 -2734 129 -2687
rect 187 -2653 287 -2637
rect 187 -2687 203 -2653
rect 271 -2687 287 -2653
rect 187 -2734 287 -2687
rect 345 -2653 445 -2637
rect 345 -2687 361 -2653
rect 429 -2687 445 -2653
rect 345 -2734 445 -2687
rect 503 -2653 603 -2637
rect 503 -2687 519 -2653
rect 587 -2687 603 -2653
rect 503 -2734 603 -2687
rect 661 -2653 761 -2637
rect 661 -2687 677 -2653
rect 745 -2687 761 -2653
rect 661 -2734 761 -2687
rect 819 -2653 919 -2637
rect 819 -2687 835 -2653
rect 903 -2687 919 -2653
rect 819 -2734 919 -2687
rect 977 -2653 1077 -2637
rect 977 -2687 993 -2653
rect 1061 -2687 1077 -2653
rect 977 -2734 1077 -2687
rect 1135 -2653 1235 -2637
rect 1135 -2687 1151 -2653
rect 1219 -2687 1235 -2653
rect 1135 -2734 1235 -2687
rect 1293 -2653 1393 -2637
rect 1293 -2687 1309 -2653
rect 1377 -2687 1393 -2653
rect 1293 -2734 1393 -2687
rect 1451 -2653 1551 -2637
rect 1451 -2687 1467 -2653
rect 1535 -2687 1551 -2653
rect 1451 -2734 1551 -2687
rect -1551 -2981 -1451 -2934
rect -1551 -3015 -1535 -2981
rect -1467 -3015 -1451 -2981
rect -1551 -3031 -1451 -3015
rect -1393 -2981 -1293 -2934
rect -1393 -3015 -1377 -2981
rect -1309 -3015 -1293 -2981
rect -1393 -3031 -1293 -3015
rect -1235 -2981 -1135 -2934
rect -1235 -3015 -1219 -2981
rect -1151 -3015 -1135 -2981
rect -1235 -3031 -1135 -3015
rect -1077 -2981 -977 -2934
rect -1077 -3015 -1061 -2981
rect -993 -3015 -977 -2981
rect -1077 -3031 -977 -3015
rect -919 -2981 -819 -2934
rect -919 -3015 -903 -2981
rect -835 -3015 -819 -2981
rect -919 -3031 -819 -3015
rect -761 -2981 -661 -2934
rect -761 -3015 -745 -2981
rect -677 -3015 -661 -2981
rect -761 -3031 -661 -3015
rect -603 -2981 -503 -2934
rect -603 -3015 -587 -2981
rect -519 -3015 -503 -2981
rect -603 -3031 -503 -3015
rect -445 -2981 -345 -2934
rect -445 -3015 -429 -2981
rect -361 -3015 -345 -2981
rect -445 -3031 -345 -3015
rect -287 -2981 -187 -2934
rect -287 -3015 -271 -2981
rect -203 -3015 -187 -2981
rect -287 -3031 -187 -3015
rect -129 -2981 -29 -2934
rect -129 -3015 -113 -2981
rect -45 -3015 -29 -2981
rect -129 -3031 -29 -3015
rect 29 -2981 129 -2934
rect 29 -3015 45 -2981
rect 113 -3015 129 -2981
rect 29 -3031 129 -3015
rect 187 -2981 287 -2934
rect 187 -3015 203 -2981
rect 271 -3015 287 -2981
rect 187 -3031 287 -3015
rect 345 -2981 445 -2934
rect 345 -3015 361 -2981
rect 429 -3015 445 -2981
rect 345 -3031 445 -3015
rect 503 -2981 603 -2934
rect 503 -3015 519 -2981
rect 587 -3015 603 -2981
rect 503 -3031 603 -3015
rect 661 -2981 761 -2934
rect 661 -3015 677 -2981
rect 745 -3015 761 -2981
rect 661 -3031 761 -3015
rect 819 -2981 919 -2934
rect 819 -3015 835 -2981
rect 903 -3015 919 -2981
rect 819 -3031 919 -3015
rect 977 -2981 1077 -2934
rect 977 -3015 993 -2981
rect 1061 -3015 1077 -2981
rect 977 -3031 1077 -3015
rect 1135 -2981 1235 -2934
rect 1135 -3015 1151 -2981
rect 1219 -3015 1235 -2981
rect 1135 -3031 1235 -3015
rect 1293 -2981 1393 -2934
rect 1293 -3015 1309 -2981
rect 1377 -3015 1393 -2981
rect 1293 -3031 1393 -3015
rect 1451 -2981 1551 -2934
rect 1451 -3015 1467 -2981
rect 1535 -3015 1551 -2981
rect 1451 -3031 1551 -3015
<< polycont >>
rect -1535 2981 -1467 3015
rect -1377 2981 -1309 3015
rect -1219 2981 -1151 3015
rect -1061 2981 -993 3015
rect -903 2981 -835 3015
rect -745 2981 -677 3015
rect -587 2981 -519 3015
rect -429 2981 -361 3015
rect -271 2981 -203 3015
rect -113 2981 -45 3015
rect 45 2981 113 3015
rect 203 2981 271 3015
rect 361 2981 429 3015
rect 519 2981 587 3015
rect 677 2981 745 3015
rect 835 2981 903 3015
rect 993 2981 1061 3015
rect 1151 2981 1219 3015
rect 1309 2981 1377 3015
rect 1467 2981 1535 3015
rect -1535 2653 -1467 2687
rect -1377 2653 -1309 2687
rect -1219 2653 -1151 2687
rect -1061 2653 -993 2687
rect -903 2653 -835 2687
rect -745 2653 -677 2687
rect -587 2653 -519 2687
rect -429 2653 -361 2687
rect -271 2653 -203 2687
rect -113 2653 -45 2687
rect 45 2653 113 2687
rect 203 2653 271 2687
rect 361 2653 429 2687
rect 519 2653 587 2687
rect 677 2653 745 2687
rect 835 2653 903 2687
rect 993 2653 1061 2687
rect 1151 2653 1219 2687
rect 1309 2653 1377 2687
rect 1467 2653 1535 2687
rect -1535 2545 -1467 2579
rect -1377 2545 -1309 2579
rect -1219 2545 -1151 2579
rect -1061 2545 -993 2579
rect -903 2545 -835 2579
rect -745 2545 -677 2579
rect -587 2545 -519 2579
rect -429 2545 -361 2579
rect -271 2545 -203 2579
rect -113 2545 -45 2579
rect 45 2545 113 2579
rect 203 2545 271 2579
rect 361 2545 429 2579
rect 519 2545 587 2579
rect 677 2545 745 2579
rect 835 2545 903 2579
rect 993 2545 1061 2579
rect 1151 2545 1219 2579
rect 1309 2545 1377 2579
rect 1467 2545 1535 2579
rect -1535 2217 -1467 2251
rect -1377 2217 -1309 2251
rect -1219 2217 -1151 2251
rect -1061 2217 -993 2251
rect -903 2217 -835 2251
rect -745 2217 -677 2251
rect -587 2217 -519 2251
rect -429 2217 -361 2251
rect -271 2217 -203 2251
rect -113 2217 -45 2251
rect 45 2217 113 2251
rect 203 2217 271 2251
rect 361 2217 429 2251
rect 519 2217 587 2251
rect 677 2217 745 2251
rect 835 2217 903 2251
rect 993 2217 1061 2251
rect 1151 2217 1219 2251
rect 1309 2217 1377 2251
rect 1467 2217 1535 2251
rect -1535 2109 -1467 2143
rect -1377 2109 -1309 2143
rect -1219 2109 -1151 2143
rect -1061 2109 -993 2143
rect -903 2109 -835 2143
rect -745 2109 -677 2143
rect -587 2109 -519 2143
rect -429 2109 -361 2143
rect -271 2109 -203 2143
rect -113 2109 -45 2143
rect 45 2109 113 2143
rect 203 2109 271 2143
rect 361 2109 429 2143
rect 519 2109 587 2143
rect 677 2109 745 2143
rect 835 2109 903 2143
rect 993 2109 1061 2143
rect 1151 2109 1219 2143
rect 1309 2109 1377 2143
rect 1467 2109 1535 2143
rect -1535 1781 -1467 1815
rect -1377 1781 -1309 1815
rect -1219 1781 -1151 1815
rect -1061 1781 -993 1815
rect -903 1781 -835 1815
rect -745 1781 -677 1815
rect -587 1781 -519 1815
rect -429 1781 -361 1815
rect -271 1781 -203 1815
rect -113 1781 -45 1815
rect 45 1781 113 1815
rect 203 1781 271 1815
rect 361 1781 429 1815
rect 519 1781 587 1815
rect 677 1781 745 1815
rect 835 1781 903 1815
rect 993 1781 1061 1815
rect 1151 1781 1219 1815
rect 1309 1781 1377 1815
rect 1467 1781 1535 1815
rect -1535 1673 -1467 1707
rect -1377 1673 -1309 1707
rect -1219 1673 -1151 1707
rect -1061 1673 -993 1707
rect -903 1673 -835 1707
rect -745 1673 -677 1707
rect -587 1673 -519 1707
rect -429 1673 -361 1707
rect -271 1673 -203 1707
rect -113 1673 -45 1707
rect 45 1673 113 1707
rect 203 1673 271 1707
rect 361 1673 429 1707
rect 519 1673 587 1707
rect 677 1673 745 1707
rect 835 1673 903 1707
rect 993 1673 1061 1707
rect 1151 1673 1219 1707
rect 1309 1673 1377 1707
rect 1467 1673 1535 1707
rect -1535 1345 -1467 1379
rect -1377 1345 -1309 1379
rect -1219 1345 -1151 1379
rect -1061 1345 -993 1379
rect -903 1345 -835 1379
rect -745 1345 -677 1379
rect -587 1345 -519 1379
rect -429 1345 -361 1379
rect -271 1345 -203 1379
rect -113 1345 -45 1379
rect 45 1345 113 1379
rect 203 1345 271 1379
rect 361 1345 429 1379
rect 519 1345 587 1379
rect 677 1345 745 1379
rect 835 1345 903 1379
rect 993 1345 1061 1379
rect 1151 1345 1219 1379
rect 1309 1345 1377 1379
rect 1467 1345 1535 1379
rect -1535 1237 -1467 1271
rect -1377 1237 -1309 1271
rect -1219 1237 -1151 1271
rect -1061 1237 -993 1271
rect -903 1237 -835 1271
rect -745 1237 -677 1271
rect -587 1237 -519 1271
rect -429 1237 -361 1271
rect -271 1237 -203 1271
rect -113 1237 -45 1271
rect 45 1237 113 1271
rect 203 1237 271 1271
rect 361 1237 429 1271
rect 519 1237 587 1271
rect 677 1237 745 1271
rect 835 1237 903 1271
rect 993 1237 1061 1271
rect 1151 1237 1219 1271
rect 1309 1237 1377 1271
rect 1467 1237 1535 1271
rect -1535 909 -1467 943
rect -1377 909 -1309 943
rect -1219 909 -1151 943
rect -1061 909 -993 943
rect -903 909 -835 943
rect -745 909 -677 943
rect -587 909 -519 943
rect -429 909 -361 943
rect -271 909 -203 943
rect -113 909 -45 943
rect 45 909 113 943
rect 203 909 271 943
rect 361 909 429 943
rect 519 909 587 943
rect 677 909 745 943
rect 835 909 903 943
rect 993 909 1061 943
rect 1151 909 1219 943
rect 1309 909 1377 943
rect 1467 909 1535 943
rect -1535 801 -1467 835
rect -1377 801 -1309 835
rect -1219 801 -1151 835
rect -1061 801 -993 835
rect -903 801 -835 835
rect -745 801 -677 835
rect -587 801 -519 835
rect -429 801 -361 835
rect -271 801 -203 835
rect -113 801 -45 835
rect 45 801 113 835
rect 203 801 271 835
rect 361 801 429 835
rect 519 801 587 835
rect 677 801 745 835
rect 835 801 903 835
rect 993 801 1061 835
rect 1151 801 1219 835
rect 1309 801 1377 835
rect 1467 801 1535 835
rect -1535 473 -1467 507
rect -1377 473 -1309 507
rect -1219 473 -1151 507
rect -1061 473 -993 507
rect -903 473 -835 507
rect -745 473 -677 507
rect -587 473 -519 507
rect -429 473 -361 507
rect -271 473 -203 507
rect -113 473 -45 507
rect 45 473 113 507
rect 203 473 271 507
rect 361 473 429 507
rect 519 473 587 507
rect 677 473 745 507
rect 835 473 903 507
rect 993 473 1061 507
rect 1151 473 1219 507
rect 1309 473 1377 507
rect 1467 473 1535 507
rect -1535 365 -1467 399
rect -1377 365 -1309 399
rect -1219 365 -1151 399
rect -1061 365 -993 399
rect -903 365 -835 399
rect -745 365 -677 399
rect -587 365 -519 399
rect -429 365 -361 399
rect -271 365 -203 399
rect -113 365 -45 399
rect 45 365 113 399
rect 203 365 271 399
rect 361 365 429 399
rect 519 365 587 399
rect 677 365 745 399
rect 835 365 903 399
rect 993 365 1061 399
rect 1151 365 1219 399
rect 1309 365 1377 399
rect 1467 365 1535 399
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect -1535 -399 -1467 -365
rect -1377 -399 -1309 -365
rect -1219 -399 -1151 -365
rect -1061 -399 -993 -365
rect -903 -399 -835 -365
rect -745 -399 -677 -365
rect -587 -399 -519 -365
rect -429 -399 -361 -365
rect -271 -399 -203 -365
rect -113 -399 -45 -365
rect 45 -399 113 -365
rect 203 -399 271 -365
rect 361 -399 429 -365
rect 519 -399 587 -365
rect 677 -399 745 -365
rect 835 -399 903 -365
rect 993 -399 1061 -365
rect 1151 -399 1219 -365
rect 1309 -399 1377 -365
rect 1467 -399 1535 -365
rect -1535 -507 -1467 -473
rect -1377 -507 -1309 -473
rect -1219 -507 -1151 -473
rect -1061 -507 -993 -473
rect -903 -507 -835 -473
rect -745 -507 -677 -473
rect -587 -507 -519 -473
rect -429 -507 -361 -473
rect -271 -507 -203 -473
rect -113 -507 -45 -473
rect 45 -507 113 -473
rect 203 -507 271 -473
rect 361 -507 429 -473
rect 519 -507 587 -473
rect 677 -507 745 -473
rect 835 -507 903 -473
rect 993 -507 1061 -473
rect 1151 -507 1219 -473
rect 1309 -507 1377 -473
rect 1467 -507 1535 -473
rect -1535 -835 -1467 -801
rect -1377 -835 -1309 -801
rect -1219 -835 -1151 -801
rect -1061 -835 -993 -801
rect -903 -835 -835 -801
rect -745 -835 -677 -801
rect -587 -835 -519 -801
rect -429 -835 -361 -801
rect -271 -835 -203 -801
rect -113 -835 -45 -801
rect 45 -835 113 -801
rect 203 -835 271 -801
rect 361 -835 429 -801
rect 519 -835 587 -801
rect 677 -835 745 -801
rect 835 -835 903 -801
rect 993 -835 1061 -801
rect 1151 -835 1219 -801
rect 1309 -835 1377 -801
rect 1467 -835 1535 -801
rect -1535 -943 -1467 -909
rect -1377 -943 -1309 -909
rect -1219 -943 -1151 -909
rect -1061 -943 -993 -909
rect -903 -943 -835 -909
rect -745 -943 -677 -909
rect -587 -943 -519 -909
rect -429 -943 -361 -909
rect -271 -943 -203 -909
rect -113 -943 -45 -909
rect 45 -943 113 -909
rect 203 -943 271 -909
rect 361 -943 429 -909
rect 519 -943 587 -909
rect 677 -943 745 -909
rect 835 -943 903 -909
rect 993 -943 1061 -909
rect 1151 -943 1219 -909
rect 1309 -943 1377 -909
rect 1467 -943 1535 -909
rect -1535 -1271 -1467 -1237
rect -1377 -1271 -1309 -1237
rect -1219 -1271 -1151 -1237
rect -1061 -1271 -993 -1237
rect -903 -1271 -835 -1237
rect -745 -1271 -677 -1237
rect -587 -1271 -519 -1237
rect -429 -1271 -361 -1237
rect -271 -1271 -203 -1237
rect -113 -1271 -45 -1237
rect 45 -1271 113 -1237
rect 203 -1271 271 -1237
rect 361 -1271 429 -1237
rect 519 -1271 587 -1237
rect 677 -1271 745 -1237
rect 835 -1271 903 -1237
rect 993 -1271 1061 -1237
rect 1151 -1271 1219 -1237
rect 1309 -1271 1377 -1237
rect 1467 -1271 1535 -1237
rect -1535 -1379 -1467 -1345
rect -1377 -1379 -1309 -1345
rect -1219 -1379 -1151 -1345
rect -1061 -1379 -993 -1345
rect -903 -1379 -835 -1345
rect -745 -1379 -677 -1345
rect -587 -1379 -519 -1345
rect -429 -1379 -361 -1345
rect -271 -1379 -203 -1345
rect -113 -1379 -45 -1345
rect 45 -1379 113 -1345
rect 203 -1379 271 -1345
rect 361 -1379 429 -1345
rect 519 -1379 587 -1345
rect 677 -1379 745 -1345
rect 835 -1379 903 -1345
rect 993 -1379 1061 -1345
rect 1151 -1379 1219 -1345
rect 1309 -1379 1377 -1345
rect 1467 -1379 1535 -1345
rect -1535 -1707 -1467 -1673
rect -1377 -1707 -1309 -1673
rect -1219 -1707 -1151 -1673
rect -1061 -1707 -993 -1673
rect -903 -1707 -835 -1673
rect -745 -1707 -677 -1673
rect -587 -1707 -519 -1673
rect -429 -1707 -361 -1673
rect -271 -1707 -203 -1673
rect -113 -1707 -45 -1673
rect 45 -1707 113 -1673
rect 203 -1707 271 -1673
rect 361 -1707 429 -1673
rect 519 -1707 587 -1673
rect 677 -1707 745 -1673
rect 835 -1707 903 -1673
rect 993 -1707 1061 -1673
rect 1151 -1707 1219 -1673
rect 1309 -1707 1377 -1673
rect 1467 -1707 1535 -1673
rect -1535 -1815 -1467 -1781
rect -1377 -1815 -1309 -1781
rect -1219 -1815 -1151 -1781
rect -1061 -1815 -993 -1781
rect -903 -1815 -835 -1781
rect -745 -1815 -677 -1781
rect -587 -1815 -519 -1781
rect -429 -1815 -361 -1781
rect -271 -1815 -203 -1781
rect -113 -1815 -45 -1781
rect 45 -1815 113 -1781
rect 203 -1815 271 -1781
rect 361 -1815 429 -1781
rect 519 -1815 587 -1781
rect 677 -1815 745 -1781
rect 835 -1815 903 -1781
rect 993 -1815 1061 -1781
rect 1151 -1815 1219 -1781
rect 1309 -1815 1377 -1781
rect 1467 -1815 1535 -1781
rect -1535 -2143 -1467 -2109
rect -1377 -2143 -1309 -2109
rect -1219 -2143 -1151 -2109
rect -1061 -2143 -993 -2109
rect -903 -2143 -835 -2109
rect -745 -2143 -677 -2109
rect -587 -2143 -519 -2109
rect -429 -2143 -361 -2109
rect -271 -2143 -203 -2109
rect -113 -2143 -45 -2109
rect 45 -2143 113 -2109
rect 203 -2143 271 -2109
rect 361 -2143 429 -2109
rect 519 -2143 587 -2109
rect 677 -2143 745 -2109
rect 835 -2143 903 -2109
rect 993 -2143 1061 -2109
rect 1151 -2143 1219 -2109
rect 1309 -2143 1377 -2109
rect 1467 -2143 1535 -2109
rect -1535 -2251 -1467 -2217
rect -1377 -2251 -1309 -2217
rect -1219 -2251 -1151 -2217
rect -1061 -2251 -993 -2217
rect -903 -2251 -835 -2217
rect -745 -2251 -677 -2217
rect -587 -2251 -519 -2217
rect -429 -2251 -361 -2217
rect -271 -2251 -203 -2217
rect -113 -2251 -45 -2217
rect 45 -2251 113 -2217
rect 203 -2251 271 -2217
rect 361 -2251 429 -2217
rect 519 -2251 587 -2217
rect 677 -2251 745 -2217
rect 835 -2251 903 -2217
rect 993 -2251 1061 -2217
rect 1151 -2251 1219 -2217
rect 1309 -2251 1377 -2217
rect 1467 -2251 1535 -2217
rect -1535 -2579 -1467 -2545
rect -1377 -2579 -1309 -2545
rect -1219 -2579 -1151 -2545
rect -1061 -2579 -993 -2545
rect -903 -2579 -835 -2545
rect -745 -2579 -677 -2545
rect -587 -2579 -519 -2545
rect -429 -2579 -361 -2545
rect -271 -2579 -203 -2545
rect -113 -2579 -45 -2545
rect 45 -2579 113 -2545
rect 203 -2579 271 -2545
rect 361 -2579 429 -2545
rect 519 -2579 587 -2545
rect 677 -2579 745 -2545
rect 835 -2579 903 -2545
rect 993 -2579 1061 -2545
rect 1151 -2579 1219 -2545
rect 1309 -2579 1377 -2545
rect 1467 -2579 1535 -2545
rect -1535 -2687 -1467 -2653
rect -1377 -2687 -1309 -2653
rect -1219 -2687 -1151 -2653
rect -1061 -2687 -993 -2653
rect -903 -2687 -835 -2653
rect -745 -2687 -677 -2653
rect -587 -2687 -519 -2653
rect -429 -2687 -361 -2653
rect -271 -2687 -203 -2653
rect -113 -2687 -45 -2653
rect 45 -2687 113 -2653
rect 203 -2687 271 -2653
rect 361 -2687 429 -2653
rect 519 -2687 587 -2653
rect 677 -2687 745 -2653
rect 835 -2687 903 -2653
rect 993 -2687 1061 -2653
rect 1151 -2687 1219 -2653
rect 1309 -2687 1377 -2653
rect 1467 -2687 1535 -2653
rect -1535 -3015 -1467 -2981
rect -1377 -3015 -1309 -2981
rect -1219 -3015 -1151 -2981
rect -1061 -3015 -993 -2981
rect -903 -3015 -835 -2981
rect -745 -3015 -677 -2981
rect -587 -3015 -519 -2981
rect -429 -3015 -361 -2981
rect -271 -3015 -203 -2981
rect -113 -3015 -45 -2981
rect 45 -3015 113 -2981
rect 203 -3015 271 -2981
rect 361 -3015 429 -2981
rect 519 -3015 587 -2981
rect 677 -3015 745 -2981
rect 835 -3015 903 -2981
rect 993 -3015 1061 -2981
rect 1151 -3015 1219 -2981
rect 1309 -3015 1377 -2981
rect 1467 -3015 1535 -2981
<< locali >>
rect -1731 3119 -1635 3153
rect 1635 3119 1731 3153
rect -1731 3057 -1697 3119
rect 1697 3057 1731 3119
rect -1551 2981 -1535 3015
rect -1467 2981 -1451 3015
rect -1393 2981 -1377 3015
rect -1309 2981 -1293 3015
rect -1235 2981 -1219 3015
rect -1151 2981 -1135 3015
rect -1077 2981 -1061 3015
rect -993 2981 -977 3015
rect -919 2981 -903 3015
rect -835 2981 -819 3015
rect -761 2981 -745 3015
rect -677 2981 -661 3015
rect -603 2981 -587 3015
rect -519 2981 -503 3015
rect -445 2981 -429 3015
rect -361 2981 -345 3015
rect -287 2981 -271 3015
rect -203 2981 -187 3015
rect -129 2981 -113 3015
rect -45 2981 -29 3015
rect 29 2981 45 3015
rect 113 2981 129 3015
rect 187 2981 203 3015
rect 271 2981 287 3015
rect 345 2981 361 3015
rect 429 2981 445 3015
rect 503 2981 519 3015
rect 587 2981 603 3015
rect 661 2981 677 3015
rect 745 2981 761 3015
rect 819 2981 835 3015
rect 903 2981 919 3015
rect 977 2981 993 3015
rect 1061 2981 1077 3015
rect 1135 2981 1151 3015
rect 1219 2981 1235 3015
rect 1293 2981 1309 3015
rect 1377 2981 1393 3015
rect 1451 2981 1467 3015
rect 1535 2981 1551 3015
rect -1597 2922 -1563 2938
rect -1597 2730 -1563 2746
rect -1439 2922 -1405 2938
rect -1439 2730 -1405 2746
rect -1281 2922 -1247 2938
rect -1281 2730 -1247 2746
rect -1123 2922 -1089 2938
rect -1123 2730 -1089 2746
rect -965 2922 -931 2938
rect -965 2730 -931 2746
rect -807 2922 -773 2938
rect -807 2730 -773 2746
rect -649 2922 -615 2938
rect -649 2730 -615 2746
rect -491 2922 -457 2938
rect -491 2730 -457 2746
rect -333 2922 -299 2938
rect -333 2730 -299 2746
rect -175 2922 -141 2938
rect -175 2730 -141 2746
rect -17 2922 17 2938
rect -17 2730 17 2746
rect 141 2922 175 2938
rect 141 2730 175 2746
rect 299 2922 333 2938
rect 299 2730 333 2746
rect 457 2922 491 2938
rect 457 2730 491 2746
rect 615 2922 649 2938
rect 615 2730 649 2746
rect 773 2922 807 2938
rect 773 2730 807 2746
rect 931 2922 965 2938
rect 931 2730 965 2746
rect 1089 2922 1123 2938
rect 1089 2730 1123 2746
rect 1247 2922 1281 2938
rect 1247 2730 1281 2746
rect 1405 2922 1439 2938
rect 1405 2730 1439 2746
rect 1563 2922 1597 2938
rect 1563 2730 1597 2746
rect -1551 2653 -1535 2687
rect -1467 2653 -1451 2687
rect -1393 2653 -1377 2687
rect -1309 2653 -1293 2687
rect -1235 2653 -1219 2687
rect -1151 2653 -1135 2687
rect -1077 2653 -1061 2687
rect -993 2653 -977 2687
rect -919 2653 -903 2687
rect -835 2653 -819 2687
rect -761 2653 -745 2687
rect -677 2653 -661 2687
rect -603 2653 -587 2687
rect -519 2653 -503 2687
rect -445 2653 -429 2687
rect -361 2653 -345 2687
rect -287 2653 -271 2687
rect -203 2653 -187 2687
rect -129 2653 -113 2687
rect -45 2653 -29 2687
rect 29 2653 45 2687
rect 113 2653 129 2687
rect 187 2653 203 2687
rect 271 2653 287 2687
rect 345 2653 361 2687
rect 429 2653 445 2687
rect 503 2653 519 2687
rect 587 2653 603 2687
rect 661 2653 677 2687
rect 745 2653 761 2687
rect 819 2653 835 2687
rect 903 2653 919 2687
rect 977 2653 993 2687
rect 1061 2653 1077 2687
rect 1135 2653 1151 2687
rect 1219 2653 1235 2687
rect 1293 2653 1309 2687
rect 1377 2653 1393 2687
rect 1451 2653 1467 2687
rect 1535 2653 1551 2687
rect -1551 2545 -1535 2579
rect -1467 2545 -1451 2579
rect -1393 2545 -1377 2579
rect -1309 2545 -1293 2579
rect -1235 2545 -1219 2579
rect -1151 2545 -1135 2579
rect -1077 2545 -1061 2579
rect -993 2545 -977 2579
rect -919 2545 -903 2579
rect -835 2545 -819 2579
rect -761 2545 -745 2579
rect -677 2545 -661 2579
rect -603 2545 -587 2579
rect -519 2545 -503 2579
rect -445 2545 -429 2579
rect -361 2545 -345 2579
rect -287 2545 -271 2579
rect -203 2545 -187 2579
rect -129 2545 -113 2579
rect -45 2545 -29 2579
rect 29 2545 45 2579
rect 113 2545 129 2579
rect 187 2545 203 2579
rect 271 2545 287 2579
rect 345 2545 361 2579
rect 429 2545 445 2579
rect 503 2545 519 2579
rect 587 2545 603 2579
rect 661 2545 677 2579
rect 745 2545 761 2579
rect 819 2545 835 2579
rect 903 2545 919 2579
rect 977 2545 993 2579
rect 1061 2545 1077 2579
rect 1135 2545 1151 2579
rect 1219 2545 1235 2579
rect 1293 2545 1309 2579
rect 1377 2545 1393 2579
rect 1451 2545 1467 2579
rect 1535 2545 1551 2579
rect -1597 2486 -1563 2502
rect -1597 2294 -1563 2310
rect -1439 2486 -1405 2502
rect -1439 2294 -1405 2310
rect -1281 2486 -1247 2502
rect -1281 2294 -1247 2310
rect -1123 2486 -1089 2502
rect -1123 2294 -1089 2310
rect -965 2486 -931 2502
rect -965 2294 -931 2310
rect -807 2486 -773 2502
rect -807 2294 -773 2310
rect -649 2486 -615 2502
rect -649 2294 -615 2310
rect -491 2486 -457 2502
rect -491 2294 -457 2310
rect -333 2486 -299 2502
rect -333 2294 -299 2310
rect -175 2486 -141 2502
rect -175 2294 -141 2310
rect -17 2486 17 2502
rect -17 2294 17 2310
rect 141 2486 175 2502
rect 141 2294 175 2310
rect 299 2486 333 2502
rect 299 2294 333 2310
rect 457 2486 491 2502
rect 457 2294 491 2310
rect 615 2486 649 2502
rect 615 2294 649 2310
rect 773 2486 807 2502
rect 773 2294 807 2310
rect 931 2486 965 2502
rect 931 2294 965 2310
rect 1089 2486 1123 2502
rect 1089 2294 1123 2310
rect 1247 2486 1281 2502
rect 1247 2294 1281 2310
rect 1405 2486 1439 2502
rect 1405 2294 1439 2310
rect 1563 2486 1597 2502
rect 1563 2294 1597 2310
rect -1551 2217 -1535 2251
rect -1467 2217 -1451 2251
rect -1393 2217 -1377 2251
rect -1309 2217 -1293 2251
rect -1235 2217 -1219 2251
rect -1151 2217 -1135 2251
rect -1077 2217 -1061 2251
rect -993 2217 -977 2251
rect -919 2217 -903 2251
rect -835 2217 -819 2251
rect -761 2217 -745 2251
rect -677 2217 -661 2251
rect -603 2217 -587 2251
rect -519 2217 -503 2251
rect -445 2217 -429 2251
rect -361 2217 -345 2251
rect -287 2217 -271 2251
rect -203 2217 -187 2251
rect -129 2217 -113 2251
rect -45 2217 -29 2251
rect 29 2217 45 2251
rect 113 2217 129 2251
rect 187 2217 203 2251
rect 271 2217 287 2251
rect 345 2217 361 2251
rect 429 2217 445 2251
rect 503 2217 519 2251
rect 587 2217 603 2251
rect 661 2217 677 2251
rect 745 2217 761 2251
rect 819 2217 835 2251
rect 903 2217 919 2251
rect 977 2217 993 2251
rect 1061 2217 1077 2251
rect 1135 2217 1151 2251
rect 1219 2217 1235 2251
rect 1293 2217 1309 2251
rect 1377 2217 1393 2251
rect 1451 2217 1467 2251
rect 1535 2217 1551 2251
rect -1551 2109 -1535 2143
rect -1467 2109 -1451 2143
rect -1393 2109 -1377 2143
rect -1309 2109 -1293 2143
rect -1235 2109 -1219 2143
rect -1151 2109 -1135 2143
rect -1077 2109 -1061 2143
rect -993 2109 -977 2143
rect -919 2109 -903 2143
rect -835 2109 -819 2143
rect -761 2109 -745 2143
rect -677 2109 -661 2143
rect -603 2109 -587 2143
rect -519 2109 -503 2143
rect -445 2109 -429 2143
rect -361 2109 -345 2143
rect -287 2109 -271 2143
rect -203 2109 -187 2143
rect -129 2109 -113 2143
rect -45 2109 -29 2143
rect 29 2109 45 2143
rect 113 2109 129 2143
rect 187 2109 203 2143
rect 271 2109 287 2143
rect 345 2109 361 2143
rect 429 2109 445 2143
rect 503 2109 519 2143
rect 587 2109 603 2143
rect 661 2109 677 2143
rect 745 2109 761 2143
rect 819 2109 835 2143
rect 903 2109 919 2143
rect 977 2109 993 2143
rect 1061 2109 1077 2143
rect 1135 2109 1151 2143
rect 1219 2109 1235 2143
rect 1293 2109 1309 2143
rect 1377 2109 1393 2143
rect 1451 2109 1467 2143
rect 1535 2109 1551 2143
rect -1597 2050 -1563 2066
rect -1597 1858 -1563 1874
rect -1439 2050 -1405 2066
rect -1439 1858 -1405 1874
rect -1281 2050 -1247 2066
rect -1281 1858 -1247 1874
rect -1123 2050 -1089 2066
rect -1123 1858 -1089 1874
rect -965 2050 -931 2066
rect -965 1858 -931 1874
rect -807 2050 -773 2066
rect -807 1858 -773 1874
rect -649 2050 -615 2066
rect -649 1858 -615 1874
rect -491 2050 -457 2066
rect -491 1858 -457 1874
rect -333 2050 -299 2066
rect -333 1858 -299 1874
rect -175 2050 -141 2066
rect -175 1858 -141 1874
rect -17 2050 17 2066
rect -17 1858 17 1874
rect 141 2050 175 2066
rect 141 1858 175 1874
rect 299 2050 333 2066
rect 299 1858 333 1874
rect 457 2050 491 2066
rect 457 1858 491 1874
rect 615 2050 649 2066
rect 615 1858 649 1874
rect 773 2050 807 2066
rect 773 1858 807 1874
rect 931 2050 965 2066
rect 931 1858 965 1874
rect 1089 2050 1123 2066
rect 1089 1858 1123 1874
rect 1247 2050 1281 2066
rect 1247 1858 1281 1874
rect 1405 2050 1439 2066
rect 1405 1858 1439 1874
rect 1563 2050 1597 2066
rect 1563 1858 1597 1874
rect -1551 1781 -1535 1815
rect -1467 1781 -1451 1815
rect -1393 1781 -1377 1815
rect -1309 1781 -1293 1815
rect -1235 1781 -1219 1815
rect -1151 1781 -1135 1815
rect -1077 1781 -1061 1815
rect -993 1781 -977 1815
rect -919 1781 -903 1815
rect -835 1781 -819 1815
rect -761 1781 -745 1815
rect -677 1781 -661 1815
rect -603 1781 -587 1815
rect -519 1781 -503 1815
rect -445 1781 -429 1815
rect -361 1781 -345 1815
rect -287 1781 -271 1815
rect -203 1781 -187 1815
rect -129 1781 -113 1815
rect -45 1781 -29 1815
rect 29 1781 45 1815
rect 113 1781 129 1815
rect 187 1781 203 1815
rect 271 1781 287 1815
rect 345 1781 361 1815
rect 429 1781 445 1815
rect 503 1781 519 1815
rect 587 1781 603 1815
rect 661 1781 677 1815
rect 745 1781 761 1815
rect 819 1781 835 1815
rect 903 1781 919 1815
rect 977 1781 993 1815
rect 1061 1781 1077 1815
rect 1135 1781 1151 1815
rect 1219 1781 1235 1815
rect 1293 1781 1309 1815
rect 1377 1781 1393 1815
rect 1451 1781 1467 1815
rect 1535 1781 1551 1815
rect -1551 1673 -1535 1707
rect -1467 1673 -1451 1707
rect -1393 1673 -1377 1707
rect -1309 1673 -1293 1707
rect -1235 1673 -1219 1707
rect -1151 1673 -1135 1707
rect -1077 1673 -1061 1707
rect -993 1673 -977 1707
rect -919 1673 -903 1707
rect -835 1673 -819 1707
rect -761 1673 -745 1707
rect -677 1673 -661 1707
rect -603 1673 -587 1707
rect -519 1673 -503 1707
rect -445 1673 -429 1707
rect -361 1673 -345 1707
rect -287 1673 -271 1707
rect -203 1673 -187 1707
rect -129 1673 -113 1707
rect -45 1673 -29 1707
rect 29 1673 45 1707
rect 113 1673 129 1707
rect 187 1673 203 1707
rect 271 1673 287 1707
rect 345 1673 361 1707
rect 429 1673 445 1707
rect 503 1673 519 1707
rect 587 1673 603 1707
rect 661 1673 677 1707
rect 745 1673 761 1707
rect 819 1673 835 1707
rect 903 1673 919 1707
rect 977 1673 993 1707
rect 1061 1673 1077 1707
rect 1135 1673 1151 1707
rect 1219 1673 1235 1707
rect 1293 1673 1309 1707
rect 1377 1673 1393 1707
rect 1451 1673 1467 1707
rect 1535 1673 1551 1707
rect -1597 1614 -1563 1630
rect -1597 1422 -1563 1438
rect -1439 1614 -1405 1630
rect -1439 1422 -1405 1438
rect -1281 1614 -1247 1630
rect -1281 1422 -1247 1438
rect -1123 1614 -1089 1630
rect -1123 1422 -1089 1438
rect -965 1614 -931 1630
rect -965 1422 -931 1438
rect -807 1614 -773 1630
rect -807 1422 -773 1438
rect -649 1614 -615 1630
rect -649 1422 -615 1438
rect -491 1614 -457 1630
rect -491 1422 -457 1438
rect -333 1614 -299 1630
rect -333 1422 -299 1438
rect -175 1614 -141 1630
rect -175 1422 -141 1438
rect -17 1614 17 1630
rect -17 1422 17 1438
rect 141 1614 175 1630
rect 141 1422 175 1438
rect 299 1614 333 1630
rect 299 1422 333 1438
rect 457 1614 491 1630
rect 457 1422 491 1438
rect 615 1614 649 1630
rect 615 1422 649 1438
rect 773 1614 807 1630
rect 773 1422 807 1438
rect 931 1614 965 1630
rect 931 1422 965 1438
rect 1089 1614 1123 1630
rect 1089 1422 1123 1438
rect 1247 1614 1281 1630
rect 1247 1422 1281 1438
rect 1405 1614 1439 1630
rect 1405 1422 1439 1438
rect 1563 1614 1597 1630
rect 1563 1422 1597 1438
rect -1551 1345 -1535 1379
rect -1467 1345 -1451 1379
rect -1393 1345 -1377 1379
rect -1309 1345 -1293 1379
rect -1235 1345 -1219 1379
rect -1151 1345 -1135 1379
rect -1077 1345 -1061 1379
rect -993 1345 -977 1379
rect -919 1345 -903 1379
rect -835 1345 -819 1379
rect -761 1345 -745 1379
rect -677 1345 -661 1379
rect -603 1345 -587 1379
rect -519 1345 -503 1379
rect -445 1345 -429 1379
rect -361 1345 -345 1379
rect -287 1345 -271 1379
rect -203 1345 -187 1379
rect -129 1345 -113 1379
rect -45 1345 -29 1379
rect 29 1345 45 1379
rect 113 1345 129 1379
rect 187 1345 203 1379
rect 271 1345 287 1379
rect 345 1345 361 1379
rect 429 1345 445 1379
rect 503 1345 519 1379
rect 587 1345 603 1379
rect 661 1345 677 1379
rect 745 1345 761 1379
rect 819 1345 835 1379
rect 903 1345 919 1379
rect 977 1345 993 1379
rect 1061 1345 1077 1379
rect 1135 1345 1151 1379
rect 1219 1345 1235 1379
rect 1293 1345 1309 1379
rect 1377 1345 1393 1379
rect 1451 1345 1467 1379
rect 1535 1345 1551 1379
rect -1551 1237 -1535 1271
rect -1467 1237 -1451 1271
rect -1393 1237 -1377 1271
rect -1309 1237 -1293 1271
rect -1235 1237 -1219 1271
rect -1151 1237 -1135 1271
rect -1077 1237 -1061 1271
rect -993 1237 -977 1271
rect -919 1237 -903 1271
rect -835 1237 -819 1271
rect -761 1237 -745 1271
rect -677 1237 -661 1271
rect -603 1237 -587 1271
rect -519 1237 -503 1271
rect -445 1237 -429 1271
rect -361 1237 -345 1271
rect -287 1237 -271 1271
rect -203 1237 -187 1271
rect -129 1237 -113 1271
rect -45 1237 -29 1271
rect 29 1237 45 1271
rect 113 1237 129 1271
rect 187 1237 203 1271
rect 271 1237 287 1271
rect 345 1237 361 1271
rect 429 1237 445 1271
rect 503 1237 519 1271
rect 587 1237 603 1271
rect 661 1237 677 1271
rect 745 1237 761 1271
rect 819 1237 835 1271
rect 903 1237 919 1271
rect 977 1237 993 1271
rect 1061 1237 1077 1271
rect 1135 1237 1151 1271
rect 1219 1237 1235 1271
rect 1293 1237 1309 1271
rect 1377 1237 1393 1271
rect 1451 1237 1467 1271
rect 1535 1237 1551 1271
rect -1597 1178 -1563 1194
rect -1597 986 -1563 1002
rect -1439 1178 -1405 1194
rect -1439 986 -1405 1002
rect -1281 1178 -1247 1194
rect -1281 986 -1247 1002
rect -1123 1178 -1089 1194
rect -1123 986 -1089 1002
rect -965 1178 -931 1194
rect -965 986 -931 1002
rect -807 1178 -773 1194
rect -807 986 -773 1002
rect -649 1178 -615 1194
rect -649 986 -615 1002
rect -491 1178 -457 1194
rect -491 986 -457 1002
rect -333 1178 -299 1194
rect -333 986 -299 1002
rect -175 1178 -141 1194
rect -175 986 -141 1002
rect -17 1178 17 1194
rect -17 986 17 1002
rect 141 1178 175 1194
rect 141 986 175 1002
rect 299 1178 333 1194
rect 299 986 333 1002
rect 457 1178 491 1194
rect 457 986 491 1002
rect 615 1178 649 1194
rect 615 986 649 1002
rect 773 1178 807 1194
rect 773 986 807 1002
rect 931 1178 965 1194
rect 931 986 965 1002
rect 1089 1178 1123 1194
rect 1089 986 1123 1002
rect 1247 1178 1281 1194
rect 1247 986 1281 1002
rect 1405 1178 1439 1194
rect 1405 986 1439 1002
rect 1563 1178 1597 1194
rect 1563 986 1597 1002
rect -1551 909 -1535 943
rect -1467 909 -1451 943
rect -1393 909 -1377 943
rect -1309 909 -1293 943
rect -1235 909 -1219 943
rect -1151 909 -1135 943
rect -1077 909 -1061 943
rect -993 909 -977 943
rect -919 909 -903 943
rect -835 909 -819 943
rect -761 909 -745 943
rect -677 909 -661 943
rect -603 909 -587 943
rect -519 909 -503 943
rect -445 909 -429 943
rect -361 909 -345 943
rect -287 909 -271 943
rect -203 909 -187 943
rect -129 909 -113 943
rect -45 909 -29 943
rect 29 909 45 943
rect 113 909 129 943
rect 187 909 203 943
rect 271 909 287 943
rect 345 909 361 943
rect 429 909 445 943
rect 503 909 519 943
rect 587 909 603 943
rect 661 909 677 943
rect 745 909 761 943
rect 819 909 835 943
rect 903 909 919 943
rect 977 909 993 943
rect 1061 909 1077 943
rect 1135 909 1151 943
rect 1219 909 1235 943
rect 1293 909 1309 943
rect 1377 909 1393 943
rect 1451 909 1467 943
rect 1535 909 1551 943
rect -1551 801 -1535 835
rect -1467 801 -1451 835
rect -1393 801 -1377 835
rect -1309 801 -1293 835
rect -1235 801 -1219 835
rect -1151 801 -1135 835
rect -1077 801 -1061 835
rect -993 801 -977 835
rect -919 801 -903 835
rect -835 801 -819 835
rect -761 801 -745 835
rect -677 801 -661 835
rect -603 801 -587 835
rect -519 801 -503 835
rect -445 801 -429 835
rect -361 801 -345 835
rect -287 801 -271 835
rect -203 801 -187 835
rect -129 801 -113 835
rect -45 801 -29 835
rect 29 801 45 835
rect 113 801 129 835
rect 187 801 203 835
rect 271 801 287 835
rect 345 801 361 835
rect 429 801 445 835
rect 503 801 519 835
rect 587 801 603 835
rect 661 801 677 835
rect 745 801 761 835
rect 819 801 835 835
rect 903 801 919 835
rect 977 801 993 835
rect 1061 801 1077 835
rect 1135 801 1151 835
rect 1219 801 1235 835
rect 1293 801 1309 835
rect 1377 801 1393 835
rect 1451 801 1467 835
rect 1535 801 1551 835
rect -1597 742 -1563 758
rect -1597 550 -1563 566
rect -1439 742 -1405 758
rect -1439 550 -1405 566
rect -1281 742 -1247 758
rect -1281 550 -1247 566
rect -1123 742 -1089 758
rect -1123 550 -1089 566
rect -965 742 -931 758
rect -965 550 -931 566
rect -807 742 -773 758
rect -807 550 -773 566
rect -649 742 -615 758
rect -649 550 -615 566
rect -491 742 -457 758
rect -491 550 -457 566
rect -333 742 -299 758
rect -333 550 -299 566
rect -175 742 -141 758
rect -175 550 -141 566
rect -17 742 17 758
rect -17 550 17 566
rect 141 742 175 758
rect 141 550 175 566
rect 299 742 333 758
rect 299 550 333 566
rect 457 742 491 758
rect 457 550 491 566
rect 615 742 649 758
rect 615 550 649 566
rect 773 742 807 758
rect 773 550 807 566
rect 931 742 965 758
rect 931 550 965 566
rect 1089 742 1123 758
rect 1089 550 1123 566
rect 1247 742 1281 758
rect 1247 550 1281 566
rect 1405 742 1439 758
rect 1405 550 1439 566
rect 1563 742 1597 758
rect 1563 550 1597 566
rect -1551 473 -1535 507
rect -1467 473 -1451 507
rect -1393 473 -1377 507
rect -1309 473 -1293 507
rect -1235 473 -1219 507
rect -1151 473 -1135 507
rect -1077 473 -1061 507
rect -993 473 -977 507
rect -919 473 -903 507
rect -835 473 -819 507
rect -761 473 -745 507
rect -677 473 -661 507
rect -603 473 -587 507
rect -519 473 -503 507
rect -445 473 -429 507
rect -361 473 -345 507
rect -287 473 -271 507
rect -203 473 -187 507
rect -129 473 -113 507
rect -45 473 -29 507
rect 29 473 45 507
rect 113 473 129 507
rect 187 473 203 507
rect 271 473 287 507
rect 345 473 361 507
rect 429 473 445 507
rect 503 473 519 507
rect 587 473 603 507
rect 661 473 677 507
rect 745 473 761 507
rect 819 473 835 507
rect 903 473 919 507
rect 977 473 993 507
rect 1061 473 1077 507
rect 1135 473 1151 507
rect 1219 473 1235 507
rect 1293 473 1309 507
rect 1377 473 1393 507
rect 1451 473 1467 507
rect 1535 473 1551 507
rect -1551 365 -1535 399
rect -1467 365 -1451 399
rect -1393 365 -1377 399
rect -1309 365 -1293 399
rect -1235 365 -1219 399
rect -1151 365 -1135 399
rect -1077 365 -1061 399
rect -993 365 -977 399
rect -919 365 -903 399
rect -835 365 -819 399
rect -761 365 -745 399
rect -677 365 -661 399
rect -603 365 -587 399
rect -519 365 -503 399
rect -445 365 -429 399
rect -361 365 -345 399
rect -287 365 -271 399
rect -203 365 -187 399
rect -129 365 -113 399
rect -45 365 -29 399
rect 29 365 45 399
rect 113 365 129 399
rect 187 365 203 399
rect 271 365 287 399
rect 345 365 361 399
rect 429 365 445 399
rect 503 365 519 399
rect 587 365 603 399
rect 661 365 677 399
rect 745 365 761 399
rect 819 365 835 399
rect 903 365 919 399
rect 977 365 993 399
rect 1061 365 1077 399
rect 1135 365 1151 399
rect 1219 365 1235 399
rect 1293 365 1309 399
rect 1377 365 1393 399
rect 1451 365 1467 399
rect 1535 365 1551 399
rect -1597 306 -1563 322
rect -1597 114 -1563 130
rect -1439 306 -1405 322
rect -1439 114 -1405 130
rect -1281 306 -1247 322
rect -1281 114 -1247 130
rect -1123 306 -1089 322
rect -1123 114 -1089 130
rect -965 306 -931 322
rect -965 114 -931 130
rect -807 306 -773 322
rect -807 114 -773 130
rect -649 306 -615 322
rect -649 114 -615 130
rect -491 306 -457 322
rect -491 114 -457 130
rect -333 306 -299 322
rect -333 114 -299 130
rect -175 306 -141 322
rect -175 114 -141 130
rect -17 306 17 322
rect -17 114 17 130
rect 141 306 175 322
rect 141 114 175 130
rect 299 306 333 322
rect 299 114 333 130
rect 457 306 491 322
rect 457 114 491 130
rect 615 306 649 322
rect 615 114 649 130
rect 773 306 807 322
rect 773 114 807 130
rect 931 306 965 322
rect 931 114 965 130
rect 1089 306 1123 322
rect 1089 114 1123 130
rect 1247 306 1281 322
rect 1247 114 1281 130
rect 1405 306 1439 322
rect 1405 114 1439 130
rect 1563 306 1597 322
rect 1563 114 1597 130
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -919 37 -903 71
rect -835 37 -819 71
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect 819 37 835 71
rect 903 37 919 71
rect 977 37 993 71
rect 1061 37 1077 71
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1451 37 1467 71
rect 1535 37 1551 71
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect -1597 -130 -1563 -114
rect -1597 -322 -1563 -306
rect -1439 -130 -1405 -114
rect -1439 -322 -1405 -306
rect -1281 -130 -1247 -114
rect -1281 -322 -1247 -306
rect -1123 -130 -1089 -114
rect -1123 -322 -1089 -306
rect -965 -130 -931 -114
rect -965 -322 -931 -306
rect -807 -130 -773 -114
rect -807 -322 -773 -306
rect -649 -130 -615 -114
rect -649 -322 -615 -306
rect -491 -130 -457 -114
rect -491 -322 -457 -306
rect -333 -130 -299 -114
rect -333 -322 -299 -306
rect -175 -130 -141 -114
rect -175 -322 -141 -306
rect -17 -130 17 -114
rect -17 -322 17 -306
rect 141 -130 175 -114
rect 141 -322 175 -306
rect 299 -130 333 -114
rect 299 -322 333 -306
rect 457 -130 491 -114
rect 457 -322 491 -306
rect 615 -130 649 -114
rect 615 -322 649 -306
rect 773 -130 807 -114
rect 773 -322 807 -306
rect 931 -130 965 -114
rect 931 -322 965 -306
rect 1089 -130 1123 -114
rect 1089 -322 1123 -306
rect 1247 -130 1281 -114
rect 1247 -322 1281 -306
rect 1405 -130 1439 -114
rect 1405 -322 1439 -306
rect 1563 -130 1597 -114
rect 1563 -322 1597 -306
rect -1551 -399 -1535 -365
rect -1467 -399 -1451 -365
rect -1393 -399 -1377 -365
rect -1309 -399 -1293 -365
rect -1235 -399 -1219 -365
rect -1151 -399 -1135 -365
rect -1077 -399 -1061 -365
rect -993 -399 -977 -365
rect -919 -399 -903 -365
rect -835 -399 -819 -365
rect -761 -399 -745 -365
rect -677 -399 -661 -365
rect -603 -399 -587 -365
rect -519 -399 -503 -365
rect -445 -399 -429 -365
rect -361 -399 -345 -365
rect -287 -399 -271 -365
rect -203 -399 -187 -365
rect -129 -399 -113 -365
rect -45 -399 -29 -365
rect 29 -399 45 -365
rect 113 -399 129 -365
rect 187 -399 203 -365
rect 271 -399 287 -365
rect 345 -399 361 -365
rect 429 -399 445 -365
rect 503 -399 519 -365
rect 587 -399 603 -365
rect 661 -399 677 -365
rect 745 -399 761 -365
rect 819 -399 835 -365
rect 903 -399 919 -365
rect 977 -399 993 -365
rect 1061 -399 1077 -365
rect 1135 -399 1151 -365
rect 1219 -399 1235 -365
rect 1293 -399 1309 -365
rect 1377 -399 1393 -365
rect 1451 -399 1467 -365
rect 1535 -399 1551 -365
rect -1551 -507 -1535 -473
rect -1467 -507 -1451 -473
rect -1393 -507 -1377 -473
rect -1309 -507 -1293 -473
rect -1235 -507 -1219 -473
rect -1151 -507 -1135 -473
rect -1077 -507 -1061 -473
rect -993 -507 -977 -473
rect -919 -507 -903 -473
rect -835 -507 -819 -473
rect -761 -507 -745 -473
rect -677 -507 -661 -473
rect -603 -507 -587 -473
rect -519 -507 -503 -473
rect -445 -507 -429 -473
rect -361 -507 -345 -473
rect -287 -507 -271 -473
rect -203 -507 -187 -473
rect -129 -507 -113 -473
rect -45 -507 -29 -473
rect 29 -507 45 -473
rect 113 -507 129 -473
rect 187 -507 203 -473
rect 271 -507 287 -473
rect 345 -507 361 -473
rect 429 -507 445 -473
rect 503 -507 519 -473
rect 587 -507 603 -473
rect 661 -507 677 -473
rect 745 -507 761 -473
rect 819 -507 835 -473
rect 903 -507 919 -473
rect 977 -507 993 -473
rect 1061 -507 1077 -473
rect 1135 -507 1151 -473
rect 1219 -507 1235 -473
rect 1293 -507 1309 -473
rect 1377 -507 1393 -473
rect 1451 -507 1467 -473
rect 1535 -507 1551 -473
rect -1597 -566 -1563 -550
rect -1597 -758 -1563 -742
rect -1439 -566 -1405 -550
rect -1439 -758 -1405 -742
rect -1281 -566 -1247 -550
rect -1281 -758 -1247 -742
rect -1123 -566 -1089 -550
rect -1123 -758 -1089 -742
rect -965 -566 -931 -550
rect -965 -758 -931 -742
rect -807 -566 -773 -550
rect -807 -758 -773 -742
rect -649 -566 -615 -550
rect -649 -758 -615 -742
rect -491 -566 -457 -550
rect -491 -758 -457 -742
rect -333 -566 -299 -550
rect -333 -758 -299 -742
rect -175 -566 -141 -550
rect -175 -758 -141 -742
rect -17 -566 17 -550
rect -17 -758 17 -742
rect 141 -566 175 -550
rect 141 -758 175 -742
rect 299 -566 333 -550
rect 299 -758 333 -742
rect 457 -566 491 -550
rect 457 -758 491 -742
rect 615 -566 649 -550
rect 615 -758 649 -742
rect 773 -566 807 -550
rect 773 -758 807 -742
rect 931 -566 965 -550
rect 931 -758 965 -742
rect 1089 -566 1123 -550
rect 1089 -758 1123 -742
rect 1247 -566 1281 -550
rect 1247 -758 1281 -742
rect 1405 -566 1439 -550
rect 1405 -758 1439 -742
rect 1563 -566 1597 -550
rect 1563 -758 1597 -742
rect -1551 -835 -1535 -801
rect -1467 -835 -1451 -801
rect -1393 -835 -1377 -801
rect -1309 -835 -1293 -801
rect -1235 -835 -1219 -801
rect -1151 -835 -1135 -801
rect -1077 -835 -1061 -801
rect -993 -835 -977 -801
rect -919 -835 -903 -801
rect -835 -835 -819 -801
rect -761 -835 -745 -801
rect -677 -835 -661 -801
rect -603 -835 -587 -801
rect -519 -835 -503 -801
rect -445 -835 -429 -801
rect -361 -835 -345 -801
rect -287 -835 -271 -801
rect -203 -835 -187 -801
rect -129 -835 -113 -801
rect -45 -835 -29 -801
rect 29 -835 45 -801
rect 113 -835 129 -801
rect 187 -835 203 -801
rect 271 -835 287 -801
rect 345 -835 361 -801
rect 429 -835 445 -801
rect 503 -835 519 -801
rect 587 -835 603 -801
rect 661 -835 677 -801
rect 745 -835 761 -801
rect 819 -835 835 -801
rect 903 -835 919 -801
rect 977 -835 993 -801
rect 1061 -835 1077 -801
rect 1135 -835 1151 -801
rect 1219 -835 1235 -801
rect 1293 -835 1309 -801
rect 1377 -835 1393 -801
rect 1451 -835 1467 -801
rect 1535 -835 1551 -801
rect -1551 -943 -1535 -909
rect -1467 -943 -1451 -909
rect -1393 -943 -1377 -909
rect -1309 -943 -1293 -909
rect -1235 -943 -1219 -909
rect -1151 -943 -1135 -909
rect -1077 -943 -1061 -909
rect -993 -943 -977 -909
rect -919 -943 -903 -909
rect -835 -943 -819 -909
rect -761 -943 -745 -909
rect -677 -943 -661 -909
rect -603 -943 -587 -909
rect -519 -943 -503 -909
rect -445 -943 -429 -909
rect -361 -943 -345 -909
rect -287 -943 -271 -909
rect -203 -943 -187 -909
rect -129 -943 -113 -909
rect -45 -943 -29 -909
rect 29 -943 45 -909
rect 113 -943 129 -909
rect 187 -943 203 -909
rect 271 -943 287 -909
rect 345 -943 361 -909
rect 429 -943 445 -909
rect 503 -943 519 -909
rect 587 -943 603 -909
rect 661 -943 677 -909
rect 745 -943 761 -909
rect 819 -943 835 -909
rect 903 -943 919 -909
rect 977 -943 993 -909
rect 1061 -943 1077 -909
rect 1135 -943 1151 -909
rect 1219 -943 1235 -909
rect 1293 -943 1309 -909
rect 1377 -943 1393 -909
rect 1451 -943 1467 -909
rect 1535 -943 1551 -909
rect -1597 -1002 -1563 -986
rect -1597 -1194 -1563 -1178
rect -1439 -1002 -1405 -986
rect -1439 -1194 -1405 -1178
rect -1281 -1002 -1247 -986
rect -1281 -1194 -1247 -1178
rect -1123 -1002 -1089 -986
rect -1123 -1194 -1089 -1178
rect -965 -1002 -931 -986
rect -965 -1194 -931 -1178
rect -807 -1002 -773 -986
rect -807 -1194 -773 -1178
rect -649 -1002 -615 -986
rect -649 -1194 -615 -1178
rect -491 -1002 -457 -986
rect -491 -1194 -457 -1178
rect -333 -1002 -299 -986
rect -333 -1194 -299 -1178
rect -175 -1002 -141 -986
rect -175 -1194 -141 -1178
rect -17 -1002 17 -986
rect -17 -1194 17 -1178
rect 141 -1002 175 -986
rect 141 -1194 175 -1178
rect 299 -1002 333 -986
rect 299 -1194 333 -1178
rect 457 -1002 491 -986
rect 457 -1194 491 -1178
rect 615 -1002 649 -986
rect 615 -1194 649 -1178
rect 773 -1002 807 -986
rect 773 -1194 807 -1178
rect 931 -1002 965 -986
rect 931 -1194 965 -1178
rect 1089 -1002 1123 -986
rect 1089 -1194 1123 -1178
rect 1247 -1002 1281 -986
rect 1247 -1194 1281 -1178
rect 1405 -1002 1439 -986
rect 1405 -1194 1439 -1178
rect 1563 -1002 1597 -986
rect 1563 -1194 1597 -1178
rect -1551 -1271 -1535 -1237
rect -1467 -1271 -1451 -1237
rect -1393 -1271 -1377 -1237
rect -1309 -1271 -1293 -1237
rect -1235 -1271 -1219 -1237
rect -1151 -1271 -1135 -1237
rect -1077 -1271 -1061 -1237
rect -993 -1271 -977 -1237
rect -919 -1271 -903 -1237
rect -835 -1271 -819 -1237
rect -761 -1271 -745 -1237
rect -677 -1271 -661 -1237
rect -603 -1271 -587 -1237
rect -519 -1271 -503 -1237
rect -445 -1271 -429 -1237
rect -361 -1271 -345 -1237
rect -287 -1271 -271 -1237
rect -203 -1271 -187 -1237
rect -129 -1271 -113 -1237
rect -45 -1271 -29 -1237
rect 29 -1271 45 -1237
rect 113 -1271 129 -1237
rect 187 -1271 203 -1237
rect 271 -1271 287 -1237
rect 345 -1271 361 -1237
rect 429 -1271 445 -1237
rect 503 -1271 519 -1237
rect 587 -1271 603 -1237
rect 661 -1271 677 -1237
rect 745 -1271 761 -1237
rect 819 -1271 835 -1237
rect 903 -1271 919 -1237
rect 977 -1271 993 -1237
rect 1061 -1271 1077 -1237
rect 1135 -1271 1151 -1237
rect 1219 -1271 1235 -1237
rect 1293 -1271 1309 -1237
rect 1377 -1271 1393 -1237
rect 1451 -1271 1467 -1237
rect 1535 -1271 1551 -1237
rect -1551 -1379 -1535 -1345
rect -1467 -1379 -1451 -1345
rect -1393 -1379 -1377 -1345
rect -1309 -1379 -1293 -1345
rect -1235 -1379 -1219 -1345
rect -1151 -1379 -1135 -1345
rect -1077 -1379 -1061 -1345
rect -993 -1379 -977 -1345
rect -919 -1379 -903 -1345
rect -835 -1379 -819 -1345
rect -761 -1379 -745 -1345
rect -677 -1379 -661 -1345
rect -603 -1379 -587 -1345
rect -519 -1379 -503 -1345
rect -445 -1379 -429 -1345
rect -361 -1379 -345 -1345
rect -287 -1379 -271 -1345
rect -203 -1379 -187 -1345
rect -129 -1379 -113 -1345
rect -45 -1379 -29 -1345
rect 29 -1379 45 -1345
rect 113 -1379 129 -1345
rect 187 -1379 203 -1345
rect 271 -1379 287 -1345
rect 345 -1379 361 -1345
rect 429 -1379 445 -1345
rect 503 -1379 519 -1345
rect 587 -1379 603 -1345
rect 661 -1379 677 -1345
rect 745 -1379 761 -1345
rect 819 -1379 835 -1345
rect 903 -1379 919 -1345
rect 977 -1379 993 -1345
rect 1061 -1379 1077 -1345
rect 1135 -1379 1151 -1345
rect 1219 -1379 1235 -1345
rect 1293 -1379 1309 -1345
rect 1377 -1379 1393 -1345
rect 1451 -1379 1467 -1345
rect 1535 -1379 1551 -1345
rect -1597 -1438 -1563 -1422
rect -1597 -1630 -1563 -1614
rect -1439 -1438 -1405 -1422
rect -1439 -1630 -1405 -1614
rect -1281 -1438 -1247 -1422
rect -1281 -1630 -1247 -1614
rect -1123 -1438 -1089 -1422
rect -1123 -1630 -1089 -1614
rect -965 -1438 -931 -1422
rect -965 -1630 -931 -1614
rect -807 -1438 -773 -1422
rect -807 -1630 -773 -1614
rect -649 -1438 -615 -1422
rect -649 -1630 -615 -1614
rect -491 -1438 -457 -1422
rect -491 -1630 -457 -1614
rect -333 -1438 -299 -1422
rect -333 -1630 -299 -1614
rect -175 -1438 -141 -1422
rect -175 -1630 -141 -1614
rect -17 -1438 17 -1422
rect -17 -1630 17 -1614
rect 141 -1438 175 -1422
rect 141 -1630 175 -1614
rect 299 -1438 333 -1422
rect 299 -1630 333 -1614
rect 457 -1438 491 -1422
rect 457 -1630 491 -1614
rect 615 -1438 649 -1422
rect 615 -1630 649 -1614
rect 773 -1438 807 -1422
rect 773 -1630 807 -1614
rect 931 -1438 965 -1422
rect 931 -1630 965 -1614
rect 1089 -1438 1123 -1422
rect 1089 -1630 1123 -1614
rect 1247 -1438 1281 -1422
rect 1247 -1630 1281 -1614
rect 1405 -1438 1439 -1422
rect 1405 -1630 1439 -1614
rect 1563 -1438 1597 -1422
rect 1563 -1630 1597 -1614
rect -1551 -1707 -1535 -1673
rect -1467 -1707 -1451 -1673
rect -1393 -1707 -1377 -1673
rect -1309 -1707 -1293 -1673
rect -1235 -1707 -1219 -1673
rect -1151 -1707 -1135 -1673
rect -1077 -1707 -1061 -1673
rect -993 -1707 -977 -1673
rect -919 -1707 -903 -1673
rect -835 -1707 -819 -1673
rect -761 -1707 -745 -1673
rect -677 -1707 -661 -1673
rect -603 -1707 -587 -1673
rect -519 -1707 -503 -1673
rect -445 -1707 -429 -1673
rect -361 -1707 -345 -1673
rect -287 -1707 -271 -1673
rect -203 -1707 -187 -1673
rect -129 -1707 -113 -1673
rect -45 -1707 -29 -1673
rect 29 -1707 45 -1673
rect 113 -1707 129 -1673
rect 187 -1707 203 -1673
rect 271 -1707 287 -1673
rect 345 -1707 361 -1673
rect 429 -1707 445 -1673
rect 503 -1707 519 -1673
rect 587 -1707 603 -1673
rect 661 -1707 677 -1673
rect 745 -1707 761 -1673
rect 819 -1707 835 -1673
rect 903 -1707 919 -1673
rect 977 -1707 993 -1673
rect 1061 -1707 1077 -1673
rect 1135 -1707 1151 -1673
rect 1219 -1707 1235 -1673
rect 1293 -1707 1309 -1673
rect 1377 -1707 1393 -1673
rect 1451 -1707 1467 -1673
rect 1535 -1707 1551 -1673
rect -1551 -1815 -1535 -1781
rect -1467 -1815 -1451 -1781
rect -1393 -1815 -1377 -1781
rect -1309 -1815 -1293 -1781
rect -1235 -1815 -1219 -1781
rect -1151 -1815 -1135 -1781
rect -1077 -1815 -1061 -1781
rect -993 -1815 -977 -1781
rect -919 -1815 -903 -1781
rect -835 -1815 -819 -1781
rect -761 -1815 -745 -1781
rect -677 -1815 -661 -1781
rect -603 -1815 -587 -1781
rect -519 -1815 -503 -1781
rect -445 -1815 -429 -1781
rect -361 -1815 -345 -1781
rect -287 -1815 -271 -1781
rect -203 -1815 -187 -1781
rect -129 -1815 -113 -1781
rect -45 -1815 -29 -1781
rect 29 -1815 45 -1781
rect 113 -1815 129 -1781
rect 187 -1815 203 -1781
rect 271 -1815 287 -1781
rect 345 -1815 361 -1781
rect 429 -1815 445 -1781
rect 503 -1815 519 -1781
rect 587 -1815 603 -1781
rect 661 -1815 677 -1781
rect 745 -1815 761 -1781
rect 819 -1815 835 -1781
rect 903 -1815 919 -1781
rect 977 -1815 993 -1781
rect 1061 -1815 1077 -1781
rect 1135 -1815 1151 -1781
rect 1219 -1815 1235 -1781
rect 1293 -1815 1309 -1781
rect 1377 -1815 1393 -1781
rect 1451 -1815 1467 -1781
rect 1535 -1815 1551 -1781
rect -1597 -1874 -1563 -1858
rect -1597 -2066 -1563 -2050
rect -1439 -1874 -1405 -1858
rect -1439 -2066 -1405 -2050
rect -1281 -1874 -1247 -1858
rect -1281 -2066 -1247 -2050
rect -1123 -1874 -1089 -1858
rect -1123 -2066 -1089 -2050
rect -965 -1874 -931 -1858
rect -965 -2066 -931 -2050
rect -807 -1874 -773 -1858
rect -807 -2066 -773 -2050
rect -649 -1874 -615 -1858
rect -649 -2066 -615 -2050
rect -491 -1874 -457 -1858
rect -491 -2066 -457 -2050
rect -333 -1874 -299 -1858
rect -333 -2066 -299 -2050
rect -175 -1874 -141 -1858
rect -175 -2066 -141 -2050
rect -17 -1874 17 -1858
rect -17 -2066 17 -2050
rect 141 -1874 175 -1858
rect 141 -2066 175 -2050
rect 299 -1874 333 -1858
rect 299 -2066 333 -2050
rect 457 -1874 491 -1858
rect 457 -2066 491 -2050
rect 615 -1874 649 -1858
rect 615 -2066 649 -2050
rect 773 -1874 807 -1858
rect 773 -2066 807 -2050
rect 931 -1874 965 -1858
rect 931 -2066 965 -2050
rect 1089 -1874 1123 -1858
rect 1089 -2066 1123 -2050
rect 1247 -1874 1281 -1858
rect 1247 -2066 1281 -2050
rect 1405 -1874 1439 -1858
rect 1405 -2066 1439 -2050
rect 1563 -1874 1597 -1858
rect 1563 -2066 1597 -2050
rect -1551 -2143 -1535 -2109
rect -1467 -2143 -1451 -2109
rect -1393 -2143 -1377 -2109
rect -1309 -2143 -1293 -2109
rect -1235 -2143 -1219 -2109
rect -1151 -2143 -1135 -2109
rect -1077 -2143 -1061 -2109
rect -993 -2143 -977 -2109
rect -919 -2143 -903 -2109
rect -835 -2143 -819 -2109
rect -761 -2143 -745 -2109
rect -677 -2143 -661 -2109
rect -603 -2143 -587 -2109
rect -519 -2143 -503 -2109
rect -445 -2143 -429 -2109
rect -361 -2143 -345 -2109
rect -287 -2143 -271 -2109
rect -203 -2143 -187 -2109
rect -129 -2143 -113 -2109
rect -45 -2143 -29 -2109
rect 29 -2143 45 -2109
rect 113 -2143 129 -2109
rect 187 -2143 203 -2109
rect 271 -2143 287 -2109
rect 345 -2143 361 -2109
rect 429 -2143 445 -2109
rect 503 -2143 519 -2109
rect 587 -2143 603 -2109
rect 661 -2143 677 -2109
rect 745 -2143 761 -2109
rect 819 -2143 835 -2109
rect 903 -2143 919 -2109
rect 977 -2143 993 -2109
rect 1061 -2143 1077 -2109
rect 1135 -2143 1151 -2109
rect 1219 -2143 1235 -2109
rect 1293 -2143 1309 -2109
rect 1377 -2143 1393 -2109
rect 1451 -2143 1467 -2109
rect 1535 -2143 1551 -2109
rect -1551 -2251 -1535 -2217
rect -1467 -2251 -1451 -2217
rect -1393 -2251 -1377 -2217
rect -1309 -2251 -1293 -2217
rect -1235 -2251 -1219 -2217
rect -1151 -2251 -1135 -2217
rect -1077 -2251 -1061 -2217
rect -993 -2251 -977 -2217
rect -919 -2251 -903 -2217
rect -835 -2251 -819 -2217
rect -761 -2251 -745 -2217
rect -677 -2251 -661 -2217
rect -603 -2251 -587 -2217
rect -519 -2251 -503 -2217
rect -445 -2251 -429 -2217
rect -361 -2251 -345 -2217
rect -287 -2251 -271 -2217
rect -203 -2251 -187 -2217
rect -129 -2251 -113 -2217
rect -45 -2251 -29 -2217
rect 29 -2251 45 -2217
rect 113 -2251 129 -2217
rect 187 -2251 203 -2217
rect 271 -2251 287 -2217
rect 345 -2251 361 -2217
rect 429 -2251 445 -2217
rect 503 -2251 519 -2217
rect 587 -2251 603 -2217
rect 661 -2251 677 -2217
rect 745 -2251 761 -2217
rect 819 -2251 835 -2217
rect 903 -2251 919 -2217
rect 977 -2251 993 -2217
rect 1061 -2251 1077 -2217
rect 1135 -2251 1151 -2217
rect 1219 -2251 1235 -2217
rect 1293 -2251 1309 -2217
rect 1377 -2251 1393 -2217
rect 1451 -2251 1467 -2217
rect 1535 -2251 1551 -2217
rect -1597 -2310 -1563 -2294
rect -1597 -2502 -1563 -2486
rect -1439 -2310 -1405 -2294
rect -1439 -2502 -1405 -2486
rect -1281 -2310 -1247 -2294
rect -1281 -2502 -1247 -2486
rect -1123 -2310 -1089 -2294
rect -1123 -2502 -1089 -2486
rect -965 -2310 -931 -2294
rect -965 -2502 -931 -2486
rect -807 -2310 -773 -2294
rect -807 -2502 -773 -2486
rect -649 -2310 -615 -2294
rect -649 -2502 -615 -2486
rect -491 -2310 -457 -2294
rect -491 -2502 -457 -2486
rect -333 -2310 -299 -2294
rect -333 -2502 -299 -2486
rect -175 -2310 -141 -2294
rect -175 -2502 -141 -2486
rect -17 -2310 17 -2294
rect -17 -2502 17 -2486
rect 141 -2310 175 -2294
rect 141 -2502 175 -2486
rect 299 -2310 333 -2294
rect 299 -2502 333 -2486
rect 457 -2310 491 -2294
rect 457 -2502 491 -2486
rect 615 -2310 649 -2294
rect 615 -2502 649 -2486
rect 773 -2310 807 -2294
rect 773 -2502 807 -2486
rect 931 -2310 965 -2294
rect 931 -2502 965 -2486
rect 1089 -2310 1123 -2294
rect 1089 -2502 1123 -2486
rect 1247 -2310 1281 -2294
rect 1247 -2502 1281 -2486
rect 1405 -2310 1439 -2294
rect 1405 -2502 1439 -2486
rect 1563 -2310 1597 -2294
rect 1563 -2502 1597 -2486
rect -1551 -2579 -1535 -2545
rect -1467 -2579 -1451 -2545
rect -1393 -2579 -1377 -2545
rect -1309 -2579 -1293 -2545
rect -1235 -2579 -1219 -2545
rect -1151 -2579 -1135 -2545
rect -1077 -2579 -1061 -2545
rect -993 -2579 -977 -2545
rect -919 -2579 -903 -2545
rect -835 -2579 -819 -2545
rect -761 -2579 -745 -2545
rect -677 -2579 -661 -2545
rect -603 -2579 -587 -2545
rect -519 -2579 -503 -2545
rect -445 -2579 -429 -2545
rect -361 -2579 -345 -2545
rect -287 -2579 -271 -2545
rect -203 -2579 -187 -2545
rect -129 -2579 -113 -2545
rect -45 -2579 -29 -2545
rect 29 -2579 45 -2545
rect 113 -2579 129 -2545
rect 187 -2579 203 -2545
rect 271 -2579 287 -2545
rect 345 -2579 361 -2545
rect 429 -2579 445 -2545
rect 503 -2579 519 -2545
rect 587 -2579 603 -2545
rect 661 -2579 677 -2545
rect 745 -2579 761 -2545
rect 819 -2579 835 -2545
rect 903 -2579 919 -2545
rect 977 -2579 993 -2545
rect 1061 -2579 1077 -2545
rect 1135 -2579 1151 -2545
rect 1219 -2579 1235 -2545
rect 1293 -2579 1309 -2545
rect 1377 -2579 1393 -2545
rect 1451 -2579 1467 -2545
rect 1535 -2579 1551 -2545
rect -1551 -2687 -1535 -2653
rect -1467 -2687 -1451 -2653
rect -1393 -2687 -1377 -2653
rect -1309 -2687 -1293 -2653
rect -1235 -2687 -1219 -2653
rect -1151 -2687 -1135 -2653
rect -1077 -2687 -1061 -2653
rect -993 -2687 -977 -2653
rect -919 -2687 -903 -2653
rect -835 -2687 -819 -2653
rect -761 -2687 -745 -2653
rect -677 -2687 -661 -2653
rect -603 -2687 -587 -2653
rect -519 -2687 -503 -2653
rect -445 -2687 -429 -2653
rect -361 -2687 -345 -2653
rect -287 -2687 -271 -2653
rect -203 -2687 -187 -2653
rect -129 -2687 -113 -2653
rect -45 -2687 -29 -2653
rect 29 -2687 45 -2653
rect 113 -2687 129 -2653
rect 187 -2687 203 -2653
rect 271 -2687 287 -2653
rect 345 -2687 361 -2653
rect 429 -2687 445 -2653
rect 503 -2687 519 -2653
rect 587 -2687 603 -2653
rect 661 -2687 677 -2653
rect 745 -2687 761 -2653
rect 819 -2687 835 -2653
rect 903 -2687 919 -2653
rect 977 -2687 993 -2653
rect 1061 -2687 1077 -2653
rect 1135 -2687 1151 -2653
rect 1219 -2687 1235 -2653
rect 1293 -2687 1309 -2653
rect 1377 -2687 1393 -2653
rect 1451 -2687 1467 -2653
rect 1535 -2687 1551 -2653
rect -1597 -2746 -1563 -2730
rect -1597 -2938 -1563 -2922
rect -1439 -2746 -1405 -2730
rect -1439 -2938 -1405 -2922
rect -1281 -2746 -1247 -2730
rect -1281 -2938 -1247 -2922
rect -1123 -2746 -1089 -2730
rect -1123 -2938 -1089 -2922
rect -965 -2746 -931 -2730
rect -965 -2938 -931 -2922
rect -807 -2746 -773 -2730
rect -807 -2938 -773 -2922
rect -649 -2746 -615 -2730
rect -649 -2938 -615 -2922
rect -491 -2746 -457 -2730
rect -491 -2938 -457 -2922
rect -333 -2746 -299 -2730
rect -333 -2938 -299 -2922
rect -175 -2746 -141 -2730
rect -175 -2938 -141 -2922
rect -17 -2746 17 -2730
rect -17 -2938 17 -2922
rect 141 -2746 175 -2730
rect 141 -2938 175 -2922
rect 299 -2746 333 -2730
rect 299 -2938 333 -2922
rect 457 -2746 491 -2730
rect 457 -2938 491 -2922
rect 615 -2746 649 -2730
rect 615 -2938 649 -2922
rect 773 -2746 807 -2730
rect 773 -2938 807 -2922
rect 931 -2746 965 -2730
rect 931 -2938 965 -2922
rect 1089 -2746 1123 -2730
rect 1089 -2938 1123 -2922
rect 1247 -2746 1281 -2730
rect 1247 -2938 1281 -2922
rect 1405 -2746 1439 -2730
rect 1405 -2938 1439 -2922
rect 1563 -2746 1597 -2730
rect 1563 -2938 1597 -2922
rect -1551 -3015 -1535 -2981
rect -1467 -3015 -1451 -2981
rect -1393 -3015 -1377 -2981
rect -1309 -3015 -1293 -2981
rect -1235 -3015 -1219 -2981
rect -1151 -3015 -1135 -2981
rect -1077 -3015 -1061 -2981
rect -993 -3015 -977 -2981
rect -919 -3015 -903 -2981
rect -835 -3015 -819 -2981
rect -761 -3015 -745 -2981
rect -677 -3015 -661 -2981
rect -603 -3015 -587 -2981
rect -519 -3015 -503 -2981
rect -445 -3015 -429 -2981
rect -361 -3015 -345 -2981
rect -287 -3015 -271 -2981
rect -203 -3015 -187 -2981
rect -129 -3015 -113 -2981
rect -45 -3015 -29 -2981
rect 29 -3015 45 -2981
rect 113 -3015 129 -2981
rect 187 -3015 203 -2981
rect 271 -3015 287 -2981
rect 345 -3015 361 -2981
rect 429 -3015 445 -2981
rect 503 -3015 519 -2981
rect 587 -3015 603 -2981
rect 661 -3015 677 -2981
rect 745 -3015 761 -2981
rect 819 -3015 835 -2981
rect 903 -3015 919 -2981
rect 977 -3015 993 -2981
rect 1061 -3015 1077 -2981
rect 1135 -3015 1151 -2981
rect 1219 -3015 1235 -2981
rect 1293 -3015 1309 -2981
rect 1377 -3015 1393 -2981
rect 1451 -3015 1467 -2981
rect 1535 -3015 1551 -2981
rect -1731 -3119 -1697 -3057
rect 1697 -3119 1731 -3057
rect -1731 -3153 -1635 -3119
rect 1635 -3153 1731 -3119
<< viali >>
rect -1535 2981 -1467 3015
rect -1377 2981 -1309 3015
rect -1219 2981 -1151 3015
rect -1061 2981 -993 3015
rect -903 2981 -835 3015
rect -745 2981 -677 3015
rect -587 2981 -519 3015
rect -429 2981 -361 3015
rect -271 2981 -203 3015
rect -113 2981 -45 3015
rect 45 2981 113 3015
rect 203 2981 271 3015
rect 361 2981 429 3015
rect 519 2981 587 3015
rect 677 2981 745 3015
rect 835 2981 903 3015
rect 993 2981 1061 3015
rect 1151 2981 1219 3015
rect 1309 2981 1377 3015
rect 1467 2981 1535 3015
rect -1597 2746 -1563 2922
rect -1439 2746 -1405 2922
rect -1281 2746 -1247 2922
rect -1123 2746 -1089 2922
rect -965 2746 -931 2922
rect -807 2746 -773 2922
rect -649 2746 -615 2922
rect -491 2746 -457 2922
rect -333 2746 -299 2922
rect -175 2746 -141 2922
rect -17 2746 17 2922
rect 141 2746 175 2922
rect 299 2746 333 2922
rect 457 2746 491 2922
rect 615 2746 649 2922
rect 773 2746 807 2922
rect 931 2746 965 2922
rect 1089 2746 1123 2922
rect 1247 2746 1281 2922
rect 1405 2746 1439 2922
rect 1563 2746 1597 2922
rect -1535 2653 -1467 2687
rect -1377 2653 -1309 2687
rect -1219 2653 -1151 2687
rect -1061 2653 -993 2687
rect -903 2653 -835 2687
rect -745 2653 -677 2687
rect -587 2653 -519 2687
rect -429 2653 -361 2687
rect -271 2653 -203 2687
rect -113 2653 -45 2687
rect 45 2653 113 2687
rect 203 2653 271 2687
rect 361 2653 429 2687
rect 519 2653 587 2687
rect 677 2653 745 2687
rect 835 2653 903 2687
rect 993 2653 1061 2687
rect 1151 2653 1219 2687
rect 1309 2653 1377 2687
rect 1467 2653 1535 2687
rect -1535 2545 -1467 2579
rect -1377 2545 -1309 2579
rect -1219 2545 -1151 2579
rect -1061 2545 -993 2579
rect -903 2545 -835 2579
rect -745 2545 -677 2579
rect -587 2545 -519 2579
rect -429 2545 -361 2579
rect -271 2545 -203 2579
rect -113 2545 -45 2579
rect 45 2545 113 2579
rect 203 2545 271 2579
rect 361 2545 429 2579
rect 519 2545 587 2579
rect 677 2545 745 2579
rect 835 2545 903 2579
rect 993 2545 1061 2579
rect 1151 2545 1219 2579
rect 1309 2545 1377 2579
rect 1467 2545 1535 2579
rect -1597 2310 -1563 2486
rect -1439 2310 -1405 2486
rect -1281 2310 -1247 2486
rect -1123 2310 -1089 2486
rect -965 2310 -931 2486
rect -807 2310 -773 2486
rect -649 2310 -615 2486
rect -491 2310 -457 2486
rect -333 2310 -299 2486
rect -175 2310 -141 2486
rect -17 2310 17 2486
rect 141 2310 175 2486
rect 299 2310 333 2486
rect 457 2310 491 2486
rect 615 2310 649 2486
rect 773 2310 807 2486
rect 931 2310 965 2486
rect 1089 2310 1123 2486
rect 1247 2310 1281 2486
rect 1405 2310 1439 2486
rect 1563 2310 1597 2486
rect -1535 2217 -1467 2251
rect -1377 2217 -1309 2251
rect -1219 2217 -1151 2251
rect -1061 2217 -993 2251
rect -903 2217 -835 2251
rect -745 2217 -677 2251
rect -587 2217 -519 2251
rect -429 2217 -361 2251
rect -271 2217 -203 2251
rect -113 2217 -45 2251
rect 45 2217 113 2251
rect 203 2217 271 2251
rect 361 2217 429 2251
rect 519 2217 587 2251
rect 677 2217 745 2251
rect 835 2217 903 2251
rect 993 2217 1061 2251
rect 1151 2217 1219 2251
rect 1309 2217 1377 2251
rect 1467 2217 1535 2251
rect -1535 2109 -1467 2143
rect -1377 2109 -1309 2143
rect -1219 2109 -1151 2143
rect -1061 2109 -993 2143
rect -903 2109 -835 2143
rect -745 2109 -677 2143
rect -587 2109 -519 2143
rect -429 2109 -361 2143
rect -271 2109 -203 2143
rect -113 2109 -45 2143
rect 45 2109 113 2143
rect 203 2109 271 2143
rect 361 2109 429 2143
rect 519 2109 587 2143
rect 677 2109 745 2143
rect 835 2109 903 2143
rect 993 2109 1061 2143
rect 1151 2109 1219 2143
rect 1309 2109 1377 2143
rect 1467 2109 1535 2143
rect -1597 1874 -1563 2050
rect -1439 1874 -1405 2050
rect -1281 1874 -1247 2050
rect -1123 1874 -1089 2050
rect -965 1874 -931 2050
rect -807 1874 -773 2050
rect -649 1874 -615 2050
rect -491 1874 -457 2050
rect -333 1874 -299 2050
rect -175 1874 -141 2050
rect -17 1874 17 2050
rect 141 1874 175 2050
rect 299 1874 333 2050
rect 457 1874 491 2050
rect 615 1874 649 2050
rect 773 1874 807 2050
rect 931 1874 965 2050
rect 1089 1874 1123 2050
rect 1247 1874 1281 2050
rect 1405 1874 1439 2050
rect 1563 1874 1597 2050
rect -1535 1781 -1467 1815
rect -1377 1781 -1309 1815
rect -1219 1781 -1151 1815
rect -1061 1781 -993 1815
rect -903 1781 -835 1815
rect -745 1781 -677 1815
rect -587 1781 -519 1815
rect -429 1781 -361 1815
rect -271 1781 -203 1815
rect -113 1781 -45 1815
rect 45 1781 113 1815
rect 203 1781 271 1815
rect 361 1781 429 1815
rect 519 1781 587 1815
rect 677 1781 745 1815
rect 835 1781 903 1815
rect 993 1781 1061 1815
rect 1151 1781 1219 1815
rect 1309 1781 1377 1815
rect 1467 1781 1535 1815
rect -1535 1673 -1467 1707
rect -1377 1673 -1309 1707
rect -1219 1673 -1151 1707
rect -1061 1673 -993 1707
rect -903 1673 -835 1707
rect -745 1673 -677 1707
rect -587 1673 -519 1707
rect -429 1673 -361 1707
rect -271 1673 -203 1707
rect -113 1673 -45 1707
rect 45 1673 113 1707
rect 203 1673 271 1707
rect 361 1673 429 1707
rect 519 1673 587 1707
rect 677 1673 745 1707
rect 835 1673 903 1707
rect 993 1673 1061 1707
rect 1151 1673 1219 1707
rect 1309 1673 1377 1707
rect 1467 1673 1535 1707
rect -1597 1438 -1563 1614
rect -1439 1438 -1405 1614
rect -1281 1438 -1247 1614
rect -1123 1438 -1089 1614
rect -965 1438 -931 1614
rect -807 1438 -773 1614
rect -649 1438 -615 1614
rect -491 1438 -457 1614
rect -333 1438 -299 1614
rect -175 1438 -141 1614
rect -17 1438 17 1614
rect 141 1438 175 1614
rect 299 1438 333 1614
rect 457 1438 491 1614
rect 615 1438 649 1614
rect 773 1438 807 1614
rect 931 1438 965 1614
rect 1089 1438 1123 1614
rect 1247 1438 1281 1614
rect 1405 1438 1439 1614
rect 1563 1438 1597 1614
rect -1535 1345 -1467 1379
rect -1377 1345 -1309 1379
rect -1219 1345 -1151 1379
rect -1061 1345 -993 1379
rect -903 1345 -835 1379
rect -745 1345 -677 1379
rect -587 1345 -519 1379
rect -429 1345 -361 1379
rect -271 1345 -203 1379
rect -113 1345 -45 1379
rect 45 1345 113 1379
rect 203 1345 271 1379
rect 361 1345 429 1379
rect 519 1345 587 1379
rect 677 1345 745 1379
rect 835 1345 903 1379
rect 993 1345 1061 1379
rect 1151 1345 1219 1379
rect 1309 1345 1377 1379
rect 1467 1345 1535 1379
rect -1535 1237 -1467 1271
rect -1377 1237 -1309 1271
rect -1219 1237 -1151 1271
rect -1061 1237 -993 1271
rect -903 1237 -835 1271
rect -745 1237 -677 1271
rect -587 1237 -519 1271
rect -429 1237 -361 1271
rect -271 1237 -203 1271
rect -113 1237 -45 1271
rect 45 1237 113 1271
rect 203 1237 271 1271
rect 361 1237 429 1271
rect 519 1237 587 1271
rect 677 1237 745 1271
rect 835 1237 903 1271
rect 993 1237 1061 1271
rect 1151 1237 1219 1271
rect 1309 1237 1377 1271
rect 1467 1237 1535 1271
rect -1597 1002 -1563 1178
rect -1439 1002 -1405 1178
rect -1281 1002 -1247 1178
rect -1123 1002 -1089 1178
rect -965 1002 -931 1178
rect -807 1002 -773 1178
rect -649 1002 -615 1178
rect -491 1002 -457 1178
rect -333 1002 -299 1178
rect -175 1002 -141 1178
rect -17 1002 17 1178
rect 141 1002 175 1178
rect 299 1002 333 1178
rect 457 1002 491 1178
rect 615 1002 649 1178
rect 773 1002 807 1178
rect 931 1002 965 1178
rect 1089 1002 1123 1178
rect 1247 1002 1281 1178
rect 1405 1002 1439 1178
rect 1563 1002 1597 1178
rect -1535 909 -1467 943
rect -1377 909 -1309 943
rect -1219 909 -1151 943
rect -1061 909 -993 943
rect -903 909 -835 943
rect -745 909 -677 943
rect -587 909 -519 943
rect -429 909 -361 943
rect -271 909 -203 943
rect -113 909 -45 943
rect 45 909 113 943
rect 203 909 271 943
rect 361 909 429 943
rect 519 909 587 943
rect 677 909 745 943
rect 835 909 903 943
rect 993 909 1061 943
rect 1151 909 1219 943
rect 1309 909 1377 943
rect 1467 909 1535 943
rect -1535 801 -1467 835
rect -1377 801 -1309 835
rect -1219 801 -1151 835
rect -1061 801 -993 835
rect -903 801 -835 835
rect -745 801 -677 835
rect -587 801 -519 835
rect -429 801 -361 835
rect -271 801 -203 835
rect -113 801 -45 835
rect 45 801 113 835
rect 203 801 271 835
rect 361 801 429 835
rect 519 801 587 835
rect 677 801 745 835
rect 835 801 903 835
rect 993 801 1061 835
rect 1151 801 1219 835
rect 1309 801 1377 835
rect 1467 801 1535 835
rect -1597 566 -1563 742
rect -1439 566 -1405 742
rect -1281 566 -1247 742
rect -1123 566 -1089 742
rect -965 566 -931 742
rect -807 566 -773 742
rect -649 566 -615 742
rect -491 566 -457 742
rect -333 566 -299 742
rect -175 566 -141 742
rect -17 566 17 742
rect 141 566 175 742
rect 299 566 333 742
rect 457 566 491 742
rect 615 566 649 742
rect 773 566 807 742
rect 931 566 965 742
rect 1089 566 1123 742
rect 1247 566 1281 742
rect 1405 566 1439 742
rect 1563 566 1597 742
rect -1535 473 -1467 507
rect -1377 473 -1309 507
rect -1219 473 -1151 507
rect -1061 473 -993 507
rect -903 473 -835 507
rect -745 473 -677 507
rect -587 473 -519 507
rect -429 473 -361 507
rect -271 473 -203 507
rect -113 473 -45 507
rect 45 473 113 507
rect 203 473 271 507
rect 361 473 429 507
rect 519 473 587 507
rect 677 473 745 507
rect 835 473 903 507
rect 993 473 1061 507
rect 1151 473 1219 507
rect 1309 473 1377 507
rect 1467 473 1535 507
rect -1535 365 -1467 399
rect -1377 365 -1309 399
rect -1219 365 -1151 399
rect -1061 365 -993 399
rect -903 365 -835 399
rect -745 365 -677 399
rect -587 365 -519 399
rect -429 365 -361 399
rect -271 365 -203 399
rect -113 365 -45 399
rect 45 365 113 399
rect 203 365 271 399
rect 361 365 429 399
rect 519 365 587 399
rect 677 365 745 399
rect 835 365 903 399
rect 993 365 1061 399
rect 1151 365 1219 399
rect 1309 365 1377 399
rect 1467 365 1535 399
rect -1597 130 -1563 306
rect -1439 130 -1405 306
rect -1281 130 -1247 306
rect -1123 130 -1089 306
rect -965 130 -931 306
rect -807 130 -773 306
rect -649 130 -615 306
rect -491 130 -457 306
rect -333 130 -299 306
rect -175 130 -141 306
rect -17 130 17 306
rect 141 130 175 306
rect 299 130 333 306
rect 457 130 491 306
rect 615 130 649 306
rect 773 130 807 306
rect 931 130 965 306
rect 1089 130 1123 306
rect 1247 130 1281 306
rect 1405 130 1439 306
rect 1563 130 1597 306
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect -1597 -306 -1563 -130
rect -1439 -306 -1405 -130
rect -1281 -306 -1247 -130
rect -1123 -306 -1089 -130
rect -965 -306 -931 -130
rect -807 -306 -773 -130
rect -649 -306 -615 -130
rect -491 -306 -457 -130
rect -333 -306 -299 -130
rect -175 -306 -141 -130
rect -17 -306 17 -130
rect 141 -306 175 -130
rect 299 -306 333 -130
rect 457 -306 491 -130
rect 615 -306 649 -130
rect 773 -306 807 -130
rect 931 -306 965 -130
rect 1089 -306 1123 -130
rect 1247 -306 1281 -130
rect 1405 -306 1439 -130
rect 1563 -306 1597 -130
rect -1535 -399 -1467 -365
rect -1377 -399 -1309 -365
rect -1219 -399 -1151 -365
rect -1061 -399 -993 -365
rect -903 -399 -835 -365
rect -745 -399 -677 -365
rect -587 -399 -519 -365
rect -429 -399 -361 -365
rect -271 -399 -203 -365
rect -113 -399 -45 -365
rect 45 -399 113 -365
rect 203 -399 271 -365
rect 361 -399 429 -365
rect 519 -399 587 -365
rect 677 -399 745 -365
rect 835 -399 903 -365
rect 993 -399 1061 -365
rect 1151 -399 1219 -365
rect 1309 -399 1377 -365
rect 1467 -399 1535 -365
rect -1535 -507 -1467 -473
rect -1377 -507 -1309 -473
rect -1219 -507 -1151 -473
rect -1061 -507 -993 -473
rect -903 -507 -835 -473
rect -745 -507 -677 -473
rect -587 -507 -519 -473
rect -429 -507 -361 -473
rect -271 -507 -203 -473
rect -113 -507 -45 -473
rect 45 -507 113 -473
rect 203 -507 271 -473
rect 361 -507 429 -473
rect 519 -507 587 -473
rect 677 -507 745 -473
rect 835 -507 903 -473
rect 993 -507 1061 -473
rect 1151 -507 1219 -473
rect 1309 -507 1377 -473
rect 1467 -507 1535 -473
rect -1597 -742 -1563 -566
rect -1439 -742 -1405 -566
rect -1281 -742 -1247 -566
rect -1123 -742 -1089 -566
rect -965 -742 -931 -566
rect -807 -742 -773 -566
rect -649 -742 -615 -566
rect -491 -742 -457 -566
rect -333 -742 -299 -566
rect -175 -742 -141 -566
rect -17 -742 17 -566
rect 141 -742 175 -566
rect 299 -742 333 -566
rect 457 -742 491 -566
rect 615 -742 649 -566
rect 773 -742 807 -566
rect 931 -742 965 -566
rect 1089 -742 1123 -566
rect 1247 -742 1281 -566
rect 1405 -742 1439 -566
rect 1563 -742 1597 -566
rect -1535 -835 -1467 -801
rect -1377 -835 -1309 -801
rect -1219 -835 -1151 -801
rect -1061 -835 -993 -801
rect -903 -835 -835 -801
rect -745 -835 -677 -801
rect -587 -835 -519 -801
rect -429 -835 -361 -801
rect -271 -835 -203 -801
rect -113 -835 -45 -801
rect 45 -835 113 -801
rect 203 -835 271 -801
rect 361 -835 429 -801
rect 519 -835 587 -801
rect 677 -835 745 -801
rect 835 -835 903 -801
rect 993 -835 1061 -801
rect 1151 -835 1219 -801
rect 1309 -835 1377 -801
rect 1467 -835 1535 -801
rect -1535 -943 -1467 -909
rect -1377 -943 -1309 -909
rect -1219 -943 -1151 -909
rect -1061 -943 -993 -909
rect -903 -943 -835 -909
rect -745 -943 -677 -909
rect -587 -943 -519 -909
rect -429 -943 -361 -909
rect -271 -943 -203 -909
rect -113 -943 -45 -909
rect 45 -943 113 -909
rect 203 -943 271 -909
rect 361 -943 429 -909
rect 519 -943 587 -909
rect 677 -943 745 -909
rect 835 -943 903 -909
rect 993 -943 1061 -909
rect 1151 -943 1219 -909
rect 1309 -943 1377 -909
rect 1467 -943 1535 -909
rect -1597 -1178 -1563 -1002
rect -1439 -1178 -1405 -1002
rect -1281 -1178 -1247 -1002
rect -1123 -1178 -1089 -1002
rect -965 -1178 -931 -1002
rect -807 -1178 -773 -1002
rect -649 -1178 -615 -1002
rect -491 -1178 -457 -1002
rect -333 -1178 -299 -1002
rect -175 -1178 -141 -1002
rect -17 -1178 17 -1002
rect 141 -1178 175 -1002
rect 299 -1178 333 -1002
rect 457 -1178 491 -1002
rect 615 -1178 649 -1002
rect 773 -1178 807 -1002
rect 931 -1178 965 -1002
rect 1089 -1178 1123 -1002
rect 1247 -1178 1281 -1002
rect 1405 -1178 1439 -1002
rect 1563 -1178 1597 -1002
rect -1535 -1271 -1467 -1237
rect -1377 -1271 -1309 -1237
rect -1219 -1271 -1151 -1237
rect -1061 -1271 -993 -1237
rect -903 -1271 -835 -1237
rect -745 -1271 -677 -1237
rect -587 -1271 -519 -1237
rect -429 -1271 -361 -1237
rect -271 -1271 -203 -1237
rect -113 -1271 -45 -1237
rect 45 -1271 113 -1237
rect 203 -1271 271 -1237
rect 361 -1271 429 -1237
rect 519 -1271 587 -1237
rect 677 -1271 745 -1237
rect 835 -1271 903 -1237
rect 993 -1271 1061 -1237
rect 1151 -1271 1219 -1237
rect 1309 -1271 1377 -1237
rect 1467 -1271 1535 -1237
rect -1535 -1379 -1467 -1345
rect -1377 -1379 -1309 -1345
rect -1219 -1379 -1151 -1345
rect -1061 -1379 -993 -1345
rect -903 -1379 -835 -1345
rect -745 -1379 -677 -1345
rect -587 -1379 -519 -1345
rect -429 -1379 -361 -1345
rect -271 -1379 -203 -1345
rect -113 -1379 -45 -1345
rect 45 -1379 113 -1345
rect 203 -1379 271 -1345
rect 361 -1379 429 -1345
rect 519 -1379 587 -1345
rect 677 -1379 745 -1345
rect 835 -1379 903 -1345
rect 993 -1379 1061 -1345
rect 1151 -1379 1219 -1345
rect 1309 -1379 1377 -1345
rect 1467 -1379 1535 -1345
rect -1597 -1614 -1563 -1438
rect -1439 -1614 -1405 -1438
rect -1281 -1614 -1247 -1438
rect -1123 -1614 -1089 -1438
rect -965 -1614 -931 -1438
rect -807 -1614 -773 -1438
rect -649 -1614 -615 -1438
rect -491 -1614 -457 -1438
rect -333 -1614 -299 -1438
rect -175 -1614 -141 -1438
rect -17 -1614 17 -1438
rect 141 -1614 175 -1438
rect 299 -1614 333 -1438
rect 457 -1614 491 -1438
rect 615 -1614 649 -1438
rect 773 -1614 807 -1438
rect 931 -1614 965 -1438
rect 1089 -1614 1123 -1438
rect 1247 -1614 1281 -1438
rect 1405 -1614 1439 -1438
rect 1563 -1614 1597 -1438
rect -1535 -1707 -1467 -1673
rect -1377 -1707 -1309 -1673
rect -1219 -1707 -1151 -1673
rect -1061 -1707 -993 -1673
rect -903 -1707 -835 -1673
rect -745 -1707 -677 -1673
rect -587 -1707 -519 -1673
rect -429 -1707 -361 -1673
rect -271 -1707 -203 -1673
rect -113 -1707 -45 -1673
rect 45 -1707 113 -1673
rect 203 -1707 271 -1673
rect 361 -1707 429 -1673
rect 519 -1707 587 -1673
rect 677 -1707 745 -1673
rect 835 -1707 903 -1673
rect 993 -1707 1061 -1673
rect 1151 -1707 1219 -1673
rect 1309 -1707 1377 -1673
rect 1467 -1707 1535 -1673
rect -1535 -1815 -1467 -1781
rect -1377 -1815 -1309 -1781
rect -1219 -1815 -1151 -1781
rect -1061 -1815 -993 -1781
rect -903 -1815 -835 -1781
rect -745 -1815 -677 -1781
rect -587 -1815 -519 -1781
rect -429 -1815 -361 -1781
rect -271 -1815 -203 -1781
rect -113 -1815 -45 -1781
rect 45 -1815 113 -1781
rect 203 -1815 271 -1781
rect 361 -1815 429 -1781
rect 519 -1815 587 -1781
rect 677 -1815 745 -1781
rect 835 -1815 903 -1781
rect 993 -1815 1061 -1781
rect 1151 -1815 1219 -1781
rect 1309 -1815 1377 -1781
rect 1467 -1815 1535 -1781
rect -1597 -2050 -1563 -1874
rect -1439 -2050 -1405 -1874
rect -1281 -2050 -1247 -1874
rect -1123 -2050 -1089 -1874
rect -965 -2050 -931 -1874
rect -807 -2050 -773 -1874
rect -649 -2050 -615 -1874
rect -491 -2050 -457 -1874
rect -333 -2050 -299 -1874
rect -175 -2050 -141 -1874
rect -17 -2050 17 -1874
rect 141 -2050 175 -1874
rect 299 -2050 333 -1874
rect 457 -2050 491 -1874
rect 615 -2050 649 -1874
rect 773 -2050 807 -1874
rect 931 -2050 965 -1874
rect 1089 -2050 1123 -1874
rect 1247 -2050 1281 -1874
rect 1405 -2050 1439 -1874
rect 1563 -2050 1597 -1874
rect -1535 -2143 -1467 -2109
rect -1377 -2143 -1309 -2109
rect -1219 -2143 -1151 -2109
rect -1061 -2143 -993 -2109
rect -903 -2143 -835 -2109
rect -745 -2143 -677 -2109
rect -587 -2143 -519 -2109
rect -429 -2143 -361 -2109
rect -271 -2143 -203 -2109
rect -113 -2143 -45 -2109
rect 45 -2143 113 -2109
rect 203 -2143 271 -2109
rect 361 -2143 429 -2109
rect 519 -2143 587 -2109
rect 677 -2143 745 -2109
rect 835 -2143 903 -2109
rect 993 -2143 1061 -2109
rect 1151 -2143 1219 -2109
rect 1309 -2143 1377 -2109
rect 1467 -2143 1535 -2109
rect -1535 -2251 -1467 -2217
rect -1377 -2251 -1309 -2217
rect -1219 -2251 -1151 -2217
rect -1061 -2251 -993 -2217
rect -903 -2251 -835 -2217
rect -745 -2251 -677 -2217
rect -587 -2251 -519 -2217
rect -429 -2251 -361 -2217
rect -271 -2251 -203 -2217
rect -113 -2251 -45 -2217
rect 45 -2251 113 -2217
rect 203 -2251 271 -2217
rect 361 -2251 429 -2217
rect 519 -2251 587 -2217
rect 677 -2251 745 -2217
rect 835 -2251 903 -2217
rect 993 -2251 1061 -2217
rect 1151 -2251 1219 -2217
rect 1309 -2251 1377 -2217
rect 1467 -2251 1535 -2217
rect -1597 -2486 -1563 -2310
rect -1439 -2486 -1405 -2310
rect -1281 -2486 -1247 -2310
rect -1123 -2486 -1089 -2310
rect -965 -2486 -931 -2310
rect -807 -2486 -773 -2310
rect -649 -2486 -615 -2310
rect -491 -2486 -457 -2310
rect -333 -2486 -299 -2310
rect -175 -2486 -141 -2310
rect -17 -2486 17 -2310
rect 141 -2486 175 -2310
rect 299 -2486 333 -2310
rect 457 -2486 491 -2310
rect 615 -2486 649 -2310
rect 773 -2486 807 -2310
rect 931 -2486 965 -2310
rect 1089 -2486 1123 -2310
rect 1247 -2486 1281 -2310
rect 1405 -2486 1439 -2310
rect 1563 -2486 1597 -2310
rect -1535 -2579 -1467 -2545
rect -1377 -2579 -1309 -2545
rect -1219 -2579 -1151 -2545
rect -1061 -2579 -993 -2545
rect -903 -2579 -835 -2545
rect -745 -2579 -677 -2545
rect -587 -2579 -519 -2545
rect -429 -2579 -361 -2545
rect -271 -2579 -203 -2545
rect -113 -2579 -45 -2545
rect 45 -2579 113 -2545
rect 203 -2579 271 -2545
rect 361 -2579 429 -2545
rect 519 -2579 587 -2545
rect 677 -2579 745 -2545
rect 835 -2579 903 -2545
rect 993 -2579 1061 -2545
rect 1151 -2579 1219 -2545
rect 1309 -2579 1377 -2545
rect 1467 -2579 1535 -2545
rect -1535 -2687 -1467 -2653
rect -1377 -2687 -1309 -2653
rect -1219 -2687 -1151 -2653
rect -1061 -2687 -993 -2653
rect -903 -2687 -835 -2653
rect -745 -2687 -677 -2653
rect -587 -2687 -519 -2653
rect -429 -2687 -361 -2653
rect -271 -2687 -203 -2653
rect -113 -2687 -45 -2653
rect 45 -2687 113 -2653
rect 203 -2687 271 -2653
rect 361 -2687 429 -2653
rect 519 -2687 587 -2653
rect 677 -2687 745 -2653
rect 835 -2687 903 -2653
rect 993 -2687 1061 -2653
rect 1151 -2687 1219 -2653
rect 1309 -2687 1377 -2653
rect 1467 -2687 1535 -2653
rect -1597 -2922 -1563 -2746
rect -1439 -2922 -1405 -2746
rect -1281 -2922 -1247 -2746
rect -1123 -2922 -1089 -2746
rect -965 -2922 -931 -2746
rect -807 -2922 -773 -2746
rect -649 -2922 -615 -2746
rect -491 -2922 -457 -2746
rect -333 -2922 -299 -2746
rect -175 -2922 -141 -2746
rect -17 -2922 17 -2746
rect 141 -2922 175 -2746
rect 299 -2922 333 -2746
rect 457 -2922 491 -2746
rect 615 -2922 649 -2746
rect 773 -2922 807 -2746
rect 931 -2922 965 -2746
rect 1089 -2922 1123 -2746
rect 1247 -2922 1281 -2746
rect 1405 -2922 1439 -2746
rect 1563 -2922 1597 -2746
rect -1535 -3015 -1467 -2981
rect -1377 -3015 -1309 -2981
rect -1219 -3015 -1151 -2981
rect -1061 -3015 -993 -2981
rect -903 -3015 -835 -2981
rect -745 -3015 -677 -2981
rect -587 -3015 -519 -2981
rect -429 -3015 -361 -2981
rect -271 -3015 -203 -2981
rect -113 -3015 -45 -2981
rect 45 -3015 113 -2981
rect 203 -3015 271 -2981
rect 361 -3015 429 -2981
rect 519 -3015 587 -2981
rect 677 -3015 745 -2981
rect 835 -3015 903 -2981
rect 993 -3015 1061 -2981
rect 1151 -3015 1219 -2981
rect 1309 -3015 1377 -2981
rect 1467 -3015 1535 -2981
<< metal1 >>
rect -1547 3015 -1455 3021
rect -1547 2981 -1535 3015
rect -1467 2981 -1455 3015
rect -1547 2975 -1455 2981
rect -1389 3015 -1297 3021
rect -1389 2981 -1377 3015
rect -1309 2981 -1297 3015
rect -1389 2975 -1297 2981
rect -1231 3015 -1139 3021
rect -1231 2981 -1219 3015
rect -1151 2981 -1139 3015
rect -1231 2975 -1139 2981
rect -1073 3015 -981 3021
rect -1073 2981 -1061 3015
rect -993 2981 -981 3015
rect -1073 2975 -981 2981
rect -915 3015 -823 3021
rect -915 2981 -903 3015
rect -835 2981 -823 3015
rect -915 2975 -823 2981
rect -757 3015 -665 3021
rect -757 2981 -745 3015
rect -677 2981 -665 3015
rect -757 2975 -665 2981
rect -599 3015 -507 3021
rect -599 2981 -587 3015
rect -519 2981 -507 3015
rect -599 2975 -507 2981
rect -441 3015 -349 3021
rect -441 2981 -429 3015
rect -361 2981 -349 3015
rect -441 2975 -349 2981
rect -283 3015 -191 3021
rect -283 2981 -271 3015
rect -203 2981 -191 3015
rect -283 2975 -191 2981
rect -125 3015 -33 3021
rect -125 2981 -113 3015
rect -45 2981 -33 3015
rect -125 2975 -33 2981
rect 33 3015 125 3021
rect 33 2981 45 3015
rect 113 2981 125 3015
rect 33 2975 125 2981
rect 191 3015 283 3021
rect 191 2981 203 3015
rect 271 2981 283 3015
rect 191 2975 283 2981
rect 349 3015 441 3021
rect 349 2981 361 3015
rect 429 2981 441 3015
rect 349 2975 441 2981
rect 507 3015 599 3021
rect 507 2981 519 3015
rect 587 2981 599 3015
rect 507 2975 599 2981
rect 665 3015 757 3021
rect 665 2981 677 3015
rect 745 2981 757 3015
rect 665 2975 757 2981
rect 823 3015 915 3021
rect 823 2981 835 3015
rect 903 2981 915 3015
rect 823 2975 915 2981
rect 981 3015 1073 3021
rect 981 2981 993 3015
rect 1061 2981 1073 3015
rect 981 2975 1073 2981
rect 1139 3015 1231 3021
rect 1139 2981 1151 3015
rect 1219 2981 1231 3015
rect 1139 2975 1231 2981
rect 1297 3015 1389 3021
rect 1297 2981 1309 3015
rect 1377 2981 1389 3015
rect 1297 2975 1389 2981
rect 1455 3015 1547 3021
rect 1455 2981 1467 3015
rect 1535 2981 1547 3015
rect 1455 2975 1547 2981
rect -1603 2922 -1557 2934
rect -1603 2746 -1597 2922
rect -1563 2746 -1557 2922
rect -1603 2734 -1557 2746
rect -1445 2922 -1399 2934
rect -1445 2746 -1439 2922
rect -1405 2746 -1399 2922
rect -1445 2734 -1399 2746
rect -1287 2922 -1241 2934
rect -1287 2746 -1281 2922
rect -1247 2746 -1241 2922
rect -1287 2734 -1241 2746
rect -1129 2922 -1083 2934
rect -1129 2746 -1123 2922
rect -1089 2746 -1083 2922
rect -1129 2734 -1083 2746
rect -971 2922 -925 2934
rect -971 2746 -965 2922
rect -931 2746 -925 2922
rect -971 2734 -925 2746
rect -813 2922 -767 2934
rect -813 2746 -807 2922
rect -773 2746 -767 2922
rect -813 2734 -767 2746
rect -655 2922 -609 2934
rect -655 2746 -649 2922
rect -615 2746 -609 2922
rect -655 2734 -609 2746
rect -497 2922 -451 2934
rect -497 2746 -491 2922
rect -457 2746 -451 2922
rect -497 2734 -451 2746
rect -339 2922 -293 2934
rect -339 2746 -333 2922
rect -299 2746 -293 2922
rect -339 2734 -293 2746
rect -181 2922 -135 2934
rect -181 2746 -175 2922
rect -141 2746 -135 2922
rect -181 2734 -135 2746
rect -23 2922 23 2934
rect -23 2746 -17 2922
rect 17 2746 23 2922
rect -23 2734 23 2746
rect 135 2922 181 2934
rect 135 2746 141 2922
rect 175 2746 181 2922
rect 135 2734 181 2746
rect 293 2922 339 2934
rect 293 2746 299 2922
rect 333 2746 339 2922
rect 293 2734 339 2746
rect 451 2922 497 2934
rect 451 2746 457 2922
rect 491 2746 497 2922
rect 451 2734 497 2746
rect 609 2922 655 2934
rect 609 2746 615 2922
rect 649 2746 655 2922
rect 609 2734 655 2746
rect 767 2922 813 2934
rect 767 2746 773 2922
rect 807 2746 813 2922
rect 767 2734 813 2746
rect 925 2922 971 2934
rect 925 2746 931 2922
rect 965 2746 971 2922
rect 925 2734 971 2746
rect 1083 2922 1129 2934
rect 1083 2746 1089 2922
rect 1123 2746 1129 2922
rect 1083 2734 1129 2746
rect 1241 2922 1287 2934
rect 1241 2746 1247 2922
rect 1281 2746 1287 2922
rect 1241 2734 1287 2746
rect 1399 2922 1445 2934
rect 1399 2746 1405 2922
rect 1439 2746 1445 2922
rect 1399 2734 1445 2746
rect 1557 2922 1603 2934
rect 1557 2746 1563 2922
rect 1597 2746 1603 2922
rect 1557 2734 1603 2746
rect -1547 2687 -1455 2693
rect -1547 2653 -1535 2687
rect -1467 2653 -1455 2687
rect -1547 2647 -1455 2653
rect -1389 2687 -1297 2693
rect -1389 2653 -1377 2687
rect -1309 2653 -1297 2687
rect -1389 2647 -1297 2653
rect -1231 2687 -1139 2693
rect -1231 2653 -1219 2687
rect -1151 2653 -1139 2687
rect -1231 2647 -1139 2653
rect -1073 2687 -981 2693
rect -1073 2653 -1061 2687
rect -993 2653 -981 2687
rect -1073 2647 -981 2653
rect -915 2687 -823 2693
rect -915 2653 -903 2687
rect -835 2653 -823 2687
rect -915 2647 -823 2653
rect -757 2687 -665 2693
rect -757 2653 -745 2687
rect -677 2653 -665 2687
rect -757 2647 -665 2653
rect -599 2687 -507 2693
rect -599 2653 -587 2687
rect -519 2653 -507 2687
rect -599 2647 -507 2653
rect -441 2687 -349 2693
rect -441 2653 -429 2687
rect -361 2653 -349 2687
rect -441 2647 -349 2653
rect -283 2687 -191 2693
rect -283 2653 -271 2687
rect -203 2653 -191 2687
rect -283 2647 -191 2653
rect -125 2687 -33 2693
rect -125 2653 -113 2687
rect -45 2653 -33 2687
rect -125 2647 -33 2653
rect 33 2687 125 2693
rect 33 2653 45 2687
rect 113 2653 125 2687
rect 33 2647 125 2653
rect 191 2687 283 2693
rect 191 2653 203 2687
rect 271 2653 283 2687
rect 191 2647 283 2653
rect 349 2687 441 2693
rect 349 2653 361 2687
rect 429 2653 441 2687
rect 349 2647 441 2653
rect 507 2687 599 2693
rect 507 2653 519 2687
rect 587 2653 599 2687
rect 507 2647 599 2653
rect 665 2687 757 2693
rect 665 2653 677 2687
rect 745 2653 757 2687
rect 665 2647 757 2653
rect 823 2687 915 2693
rect 823 2653 835 2687
rect 903 2653 915 2687
rect 823 2647 915 2653
rect 981 2687 1073 2693
rect 981 2653 993 2687
rect 1061 2653 1073 2687
rect 981 2647 1073 2653
rect 1139 2687 1231 2693
rect 1139 2653 1151 2687
rect 1219 2653 1231 2687
rect 1139 2647 1231 2653
rect 1297 2687 1389 2693
rect 1297 2653 1309 2687
rect 1377 2653 1389 2687
rect 1297 2647 1389 2653
rect 1455 2687 1547 2693
rect 1455 2653 1467 2687
rect 1535 2653 1547 2687
rect 1455 2647 1547 2653
rect -1547 2579 -1455 2585
rect -1547 2545 -1535 2579
rect -1467 2545 -1455 2579
rect -1547 2539 -1455 2545
rect -1389 2579 -1297 2585
rect -1389 2545 -1377 2579
rect -1309 2545 -1297 2579
rect -1389 2539 -1297 2545
rect -1231 2579 -1139 2585
rect -1231 2545 -1219 2579
rect -1151 2545 -1139 2579
rect -1231 2539 -1139 2545
rect -1073 2579 -981 2585
rect -1073 2545 -1061 2579
rect -993 2545 -981 2579
rect -1073 2539 -981 2545
rect -915 2579 -823 2585
rect -915 2545 -903 2579
rect -835 2545 -823 2579
rect -915 2539 -823 2545
rect -757 2579 -665 2585
rect -757 2545 -745 2579
rect -677 2545 -665 2579
rect -757 2539 -665 2545
rect -599 2579 -507 2585
rect -599 2545 -587 2579
rect -519 2545 -507 2579
rect -599 2539 -507 2545
rect -441 2579 -349 2585
rect -441 2545 -429 2579
rect -361 2545 -349 2579
rect -441 2539 -349 2545
rect -283 2579 -191 2585
rect -283 2545 -271 2579
rect -203 2545 -191 2579
rect -283 2539 -191 2545
rect -125 2579 -33 2585
rect -125 2545 -113 2579
rect -45 2545 -33 2579
rect -125 2539 -33 2545
rect 33 2579 125 2585
rect 33 2545 45 2579
rect 113 2545 125 2579
rect 33 2539 125 2545
rect 191 2579 283 2585
rect 191 2545 203 2579
rect 271 2545 283 2579
rect 191 2539 283 2545
rect 349 2579 441 2585
rect 349 2545 361 2579
rect 429 2545 441 2579
rect 349 2539 441 2545
rect 507 2579 599 2585
rect 507 2545 519 2579
rect 587 2545 599 2579
rect 507 2539 599 2545
rect 665 2579 757 2585
rect 665 2545 677 2579
rect 745 2545 757 2579
rect 665 2539 757 2545
rect 823 2579 915 2585
rect 823 2545 835 2579
rect 903 2545 915 2579
rect 823 2539 915 2545
rect 981 2579 1073 2585
rect 981 2545 993 2579
rect 1061 2545 1073 2579
rect 981 2539 1073 2545
rect 1139 2579 1231 2585
rect 1139 2545 1151 2579
rect 1219 2545 1231 2579
rect 1139 2539 1231 2545
rect 1297 2579 1389 2585
rect 1297 2545 1309 2579
rect 1377 2545 1389 2579
rect 1297 2539 1389 2545
rect 1455 2579 1547 2585
rect 1455 2545 1467 2579
rect 1535 2545 1547 2579
rect 1455 2539 1547 2545
rect -1603 2486 -1557 2498
rect -1603 2310 -1597 2486
rect -1563 2310 -1557 2486
rect -1603 2298 -1557 2310
rect -1445 2486 -1399 2498
rect -1445 2310 -1439 2486
rect -1405 2310 -1399 2486
rect -1445 2298 -1399 2310
rect -1287 2486 -1241 2498
rect -1287 2310 -1281 2486
rect -1247 2310 -1241 2486
rect -1287 2298 -1241 2310
rect -1129 2486 -1083 2498
rect -1129 2310 -1123 2486
rect -1089 2310 -1083 2486
rect -1129 2298 -1083 2310
rect -971 2486 -925 2498
rect -971 2310 -965 2486
rect -931 2310 -925 2486
rect -971 2298 -925 2310
rect -813 2486 -767 2498
rect -813 2310 -807 2486
rect -773 2310 -767 2486
rect -813 2298 -767 2310
rect -655 2486 -609 2498
rect -655 2310 -649 2486
rect -615 2310 -609 2486
rect -655 2298 -609 2310
rect -497 2486 -451 2498
rect -497 2310 -491 2486
rect -457 2310 -451 2486
rect -497 2298 -451 2310
rect -339 2486 -293 2498
rect -339 2310 -333 2486
rect -299 2310 -293 2486
rect -339 2298 -293 2310
rect -181 2486 -135 2498
rect -181 2310 -175 2486
rect -141 2310 -135 2486
rect -181 2298 -135 2310
rect -23 2486 23 2498
rect -23 2310 -17 2486
rect 17 2310 23 2486
rect -23 2298 23 2310
rect 135 2486 181 2498
rect 135 2310 141 2486
rect 175 2310 181 2486
rect 135 2298 181 2310
rect 293 2486 339 2498
rect 293 2310 299 2486
rect 333 2310 339 2486
rect 293 2298 339 2310
rect 451 2486 497 2498
rect 451 2310 457 2486
rect 491 2310 497 2486
rect 451 2298 497 2310
rect 609 2486 655 2498
rect 609 2310 615 2486
rect 649 2310 655 2486
rect 609 2298 655 2310
rect 767 2486 813 2498
rect 767 2310 773 2486
rect 807 2310 813 2486
rect 767 2298 813 2310
rect 925 2486 971 2498
rect 925 2310 931 2486
rect 965 2310 971 2486
rect 925 2298 971 2310
rect 1083 2486 1129 2498
rect 1083 2310 1089 2486
rect 1123 2310 1129 2486
rect 1083 2298 1129 2310
rect 1241 2486 1287 2498
rect 1241 2310 1247 2486
rect 1281 2310 1287 2486
rect 1241 2298 1287 2310
rect 1399 2486 1445 2498
rect 1399 2310 1405 2486
rect 1439 2310 1445 2486
rect 1399 2298 1445 2310
rect 1557 2486 1603 2498
rect 1557 2310 1563 2486
rect 1597 2310 1603 2486
rect 1557 2298 1603 2310
rect -1547 2251 -1455 2257
rect -1547 2217 -1535 2251
rect -1467 2217 -1455 2251
rect -1547 2211 -1455 2217
rect -1389 2251 -1297 2257
rect -1389 2217 -1377 2251
rect -1309 2217 -1297 2251
rect -1389 2211 -1297 2217
rect -1231 2251 -1139 2257
rect -1231 2217 -1219 2251
rect -1151 2217 -1139 2251
rect -1231 2211 -1139 2217
rect -1073 2251 -981 2257
rect -1073 2217 -1061 2251
rect -993 2217 -981 2251
rect -1073 2211 -981 2217
rect -915 2251 -823 2257
rect -915 2217 -903 2251
rect -835 2217 -823 2251
rect -915 2211 -823 2217
rect -757 2251 -665 2257
rect -757 2217 -745 2251
rect -677 2217 -665 2251
rect -757 2211 -665 2217
rect -599 2251 -507 2257
rect -599 2217 -587 2251
rect -519 2217 -507 2251
rect -599 2211 -507 2217
rect -441 2251 -349 2257
rect -441 2217 -429 2251
rect -361 2217 -349 2251
rect -441 2211 -349 2217
rect -283 2251 -191 2257
rect -283 2217 -271 2251
rect -203 2217 -191 2251
rect -283 2211 -191 2217
rect -125 2251 -33 2257
rect -125 2217 -113 2251
rect -45 2217 -33 2251
rect -125 2211 -33 2217
rect 33 2251 125 2257
rect 33 2217 45 2251
rect 113 2217 125 2251
rect 33 2211 125 2217
rect 191 2251 283 2257
rect 191 2217 203 2251
rect 271 2217 283 2251
rect 191 2211 283 2217
rect 349 2251 441 2257
rect 349 2217 361 2251
rect 429 2217 441 2251
rect 349 2211 441 2217
rect 507 2251 599 2257
rect 507 2217 519 2251
rect 587 2217 599 2251
rect 507 2211 599 2217
rect 665 2251 757 2257
rect 665 2217 677 2251
rect 745 2217 757 2251
rect 665 2211 757 2217
rect 823 2251 915 2257
rect 823 2217 835 2251
rect 903 2217 915 2251
rect 823 2211 915 2217
rect 981 2251 1073 2257
rect 981 2217 993 2251
rect 1061 2217 1073 2251
rect 981 2211 1073 2217
rect 1139 2251 1231 2257
rect 1139 2217 1151 2251
rect 1219 2217 1231 2251
rect 1139 2211 1231 2217
rect 1297 2251 1389 2257
rect 1297 2217 1309 2251
rect 1377 2217 1389 2251
rect 1297 2211 1389 2217
rect 1455 2251 1547 2257
rect 1455 2217 1467 2251
rect 1535 2217 1547 2251
rect 1455 2211 1547 2217
rect -1547 2143 -1455 2149
rect -1547 2109 -1535 2143
rect -1467 2109 -1455 2143
rect -1547 2103 -1455 2109
rect -1389 2143 -1297 2149
rect -1389 2109 -1377 2143
rect -1309 2109 -1297 2143
rect -1389 2103 -1297 2109
rect -1231 2143 -1139 2149
rect -1231 2109 -1219 2143
rect -1151 2109 -1139 2143
rect -1231 2103 -1139 2109
rect -1073 2143 -981 2149
rect -1073 2109 -1061 2143
rect -993 2109 -981 2143
rect -1073 2103 -981 2109
rect -915 2143 -823 2149
rect -915 2109 -903 2143
rect -835 2109 -823 2143
rect -915 2103 -823 2109
rect -757 2143 -665 2149
rect -757 2109 -745 2143
rect -677 2109 -665 2143
rect -757 2103 -665 2109
rect -599 2143 -507 2149
rect -599 2109 -587 2143
rect -519 2109 -507 2143
rect -599 2103 -507 2109
rect -441 2143 -349 2149
rect -441 2109 -429 2143
rect -361 2109 -349 2143
rect -441 2103 -349 2109
rect -283 2143 -191 2149
rect -283 2109 -271 2143
rect -203 2109 -191 2143
rect -283 2103 -191 2109
rect -125 2143 -33 2149
rect -125 2109 -113 2143
rect -45 2109 -33 2143
rect -125 2103 -33 2109
rect 33 2143 125 2149
rect 33 2109 45 2143
rect 113 2109 125 2143
rect 33 2103 125 2109
rect 191 2143 283 2149
rect 191 2109 203 2143
rect 271 2109 283 2143
rect 191 2103 283 2109
rect 349 2143 441 2149
rect 349 2109 361 2143
rect 429 2109 441 2143
rect 349 2103 441 2109
rect 507 2143 599 2149
rect 507 2109 519 2143
rect 587 2109 599 2143
rect 507 2103 599 2109
rect 665 2143 757 2149
rect 665 2109 677 2143
rect 745 2109 757 2143
rect 665 2103 757 2109
rect 823 2143 915 2149
rect 823 2109 835 2143
rect 903 2109 915 2143
rect 823 2103 915 2109
rect 981 2143 1073 2149
rect 981 2109 993 2143
rect 1061 2109 1073 2143
rect 981 2103 1073 2109
rect 1139 2143 1231 2149
rect 1139 2109 1151 2143
rect 1219 2109 1231 2143
rect 1139 2103 1231 2109
rect 1297 2143 1389 2149
rect 1297 2109 1309 2143
rect 1377 2109 1389 2143
rect 1297 2103 1389 2109
rect 1455 2143 1547 2149
rect 1455 2109 1467 2143
rect 1535 2109 1547 2143
rect 1455 2103 1547 2109
rect -1603 2050 -1557 2062
rect -1603 1874 -1597 2050
rect -1563 1874 -1557 2050
rect -1603 1862 -1557 1874
rect -1445 2050 -1399 2062
rect -1445 1874 -1439 2050
rect -1405 1874 -1399 2050
rect -1445 1862 -1399 1874
rect -1287 2050 -1241 2062
rect -1287 1874 -1281 2050
rect -1247 1874 -1241 2050
rect -1287 1862 -1241 1874
rect -1129 2050 -1083 2062
rect -1129 1874 -1123 2050
rect -1089 1874 -1083 2050
rect -1129 1862 -1083 1874
rect -971 2050 -925 2062
rect -971 1874 -965 2050
rect -931 1874 -925 2050
rect -971 1862 -925 1874
rect -813 2050 -767 2062
rect -813 1874 -807 2050
rect -773 1874 -767 2050
rect -813 1862 -767 1874
rect -655 2050 -609 2062
rect -655 1874 -649 2050
rect -615 1874 -609 2050
rect -655 1862 -609 1874
rect -497 2050 -451 2062
rect -497 1874 -491 2050
rect -457 1874 -451 2050
rect -497 1862 -451 1874
rect -339 2050 -293 2062
rect -339 1874 -333 2050
rect -299 1874 -293 2050
rect -339 1862 -293 1874
rect -181 2050 -135 2062
rect -181 1874 -175 2050
rect -141 1874 -135 2050
rect -181 1862 -135 1874
rect -23 2050 23 2062
rect -23 1874 -17 2050
rect 17 1874 23 2050
rect -23 1862 23 1874
rect 135 2050 181 2062
rect 135 1874 141 2050
rect 175 1874 181 2050
rect 135 1862 181 1874
rect 293 2050 339 2062
rect 293 1874 299 2050
rect 333 1874 339 2050
rect 293 1862 339 1874
rect 451 2050 497 2062
rect 451 1874 457 2050
rect 491 1874 497 2050
rect 451 1862 497 1874
rect 609 2050 655 2062
rect 609 1874 615 2050
rect 649 1874 655 2050
rect 609 1862 655 1874
rect 767 2050 813 2062
rect 767 1874 773 2050
rect 807 1874 813 2050
rect 767 1862 813 1874
rect 925 2050 971 2062
rect 925 1874 931 2050
rect 965 1874 971 2050
rect 925 1862 971 1874
rect 1083 2050 1129 2062
rect 1083 1874 1089 2050
rect 1123 1874 1129 2050
rect 1083 1862 1129 1874
rect 1241 2050 1287 2062
rect 1241 1874 1247 2050
rect 1281 1874 1287 2050
rect 1241 1862 1287 1874
rect 1399 2050 1445 2062
rect 1399 1874 1405 2050
rect 1439 1874 1445 2050
rect 1399 1862 1445 1874
rect 1557 2050 1603 2062
rect 1557 1874 1563 2050
rect 1597 1874 1603 2050
rect 1557 1862 1603 1874
rect -1547 1815 -1455 1821
rect -1547 1781 -1535 1815
rect -1467 1781 -1455 1815
rect -1547 1775 -1455 1781
rect -1389 1815 -1297 1821
rect -1389 1781 -1377 1815
rect -1309 1781 -1297 1815
rect -1389 1775 -1297 1781
rect -1231 1815 -1139 1821
rect -1231 1781 -1219 1815
rect -1151 1781 -1139 1815
rect -1231 1775 -1139 1781
rect -1073 1815 -981 1821
rect -1073 1781 -1061 1815
rect -993 1781 -981 1815
rect -1073 1775 -981 1781
rect -915 1815 -823 1821
rect -915 1781 -903 1815
rect -835 1781 -823 1815
rect -915 1775 -823 1781
rect -757 1815 -665 1821
rect -757 1781 -745 1815
rect -677 1781 -665 1815
rect -757 1775 -665 1781
rect -599 1815 -507 1821
rect -599 1781 -587 1815
rect -519 1781 -507 1815
rect -599 1775 -507 1781
rect -441 1815 -349 1821
rect -441 1781 -429 1815
rect -361 1781 -349 1815
rect -441 1775 -349 1781
rect -283 1815 -191 1821
rect -283 1781 -271 1815
rect -203 1781 -191 1815
rect -283 1775 -191 1781
rect -125 1815 -33 1821
rect -125 1781 -113 1815
rect -45 1781 -33 1815
rect -125 1775 -33 1781
rect 33 1815 125 1821
rect 33 1781 45 1815
rect 113 1781 125 1815
rect 33 1775 125 1781
rect 191 1815 283 1821
rect 191 1781 203 1815
rect 271 1781 283 1815
rect 191 1775 283 1781
rect 349 1815 441 1821
rect 349 1781 361 1815
rect 429 1781 441 1815
rect 349 1775 441 1781
rect 507 1815 599 1821
rect 507 1781 519 1815
rect 587 1781 599 1815
rect 507 1775 599 1781
rect 665 1815 757 1821
rect 665 1781 677 1815
rect 745 1781 757 1815
rect 665 1775 757 1781
rect 823 1815 915 1821
rect 823 1781 835 1815
rect 903 1781 915 1815
rect 823 1775 915 1781
rect 981 1815 1073 1821
rect 981 1781 993 1815
rect 1061 1781 1073 1815
rect 981 1775 1073 1781
rect 1139 1815 1231 1821
rect 1139 1781 1151 1815
rect 1219 1781 1231 1815
rect 1139 1775 1231 1781
rect 1297 1815 1389 1821
rect 1297 1781 1309 1815
rect 1377 1781 1389 1815
rect 1297 1775 1389 1781
rect 1455 1815 1547 1821
rect 1455 1781 1467 1815
rect 1535 1781 1547 1815
rect 1455 1775 1547 1781
rect -1547 1707 -1455 1713
rect -1547 1673 -1535 1707
rect -1467 1673 -1455 1707
rect -1547 1667 -1455 1673
rect -1389 1707 -1297 1713
rect -1389 1673 -1377 1707
rect -1309 1673 -1297 1707
rect -1389 1667 -1297 1673
rect -1231 1707 -1139 1713
rect -1231 1673 -1219 1707
rect -1151 1673 -1139 1707
rect -1231 1667 -1139 1673
rect -1073 1707 -981 1713
rect -1073 1673 -1061 1707
rect -993 1673 -981 1707
rect -1073 1667 -981 1673
rect -915 1707 -823 1713
rect -915 1673 -903 1707
rect -835 1673 -823 1707
rect -915 1667 -823 1673
rect -757 1707 -665 1713
rect -757 1673 -745 1707
rect -677 1673 -665 1707
rect -757 1667 -665 1673
rect -599 1707 -507 1713
rect -599 1673 -587 1707
rect -519 1673 -507 1707
rect -599 1667 -507 1673
rect -441 1707 -349 1713
rect -441 1673 -429 1707
rect -361 1673 -349 1707
rect -441 1667 -349 1673
rect -283 1707 -191 1713
rect -283 1673 -271 1707
rect -203 1673 -191 1707
rect -283 1667 -191 1673
rect -125 1707 -33 1713
rect -125 1673 -113 1707
rect -45 1673 -33 1707
rect -125 1667 -33 1673
rect 33 1707 125 1713
rect 33 1673 45 1707
rect 113 1673 125 1707
rect 33 1667 125 1673
rect 191 1707 283 1713
rect 191 1673 203 1707
rect 271 1673 283 1707
rect 191 1667 283 1673
rect 349 1707 441 1713
rect 349 1673 361 1707
rect 429 1673 441 1707
rect 349 1667 441 1673
rect 507 1707 599 1713
rect 507 1673 519 1707
rect 587 1673 599 1707
rect 507 1667 599 1673
rect 665 1707 757 1713
rect 665 1673 677 1707
rect 745 1673 757 1707
rect 665 1667 757 1673
rect 823 1707 915 1713
rect 823 1673 835 1707
rect 903 1673 915 1707
rect 823 1667 915 1673
rect 981 1707 1073 1713
rect 981 1673 993 1707
rect 1061 1673 1073 1707
rect 981 1667 1073 1673
rect 1139 1707 1231 1713
rect 1139 1673 1151 1707
rect 1219 1673 1231 1707
rect 1139 1667 1231 1673
rect 1297 1707 1389 1713
rect 1297 1673 1309 1707
rect 1377 1673 1389 1707
rect 1297 1667 1389 1673
rect 1455 1707 1547 1713
rect 1455 1673 1467 1707
rect 1535 1673 1547 1707
rect 1455 1667 1547 1673
rect -1603 1614 -1557 1626
rect -1603 1438 -1597 1614
rect -1563 1438 -1557 1614
rect -1603 1426 -1557 1438
rect -1445 1614 -1399 1626
rect -1445 1438 -1439 1614
rect -1405 1438 -1399 1614
rect -1445 1426 -1399 1438
rect -1287 1614 -1241 1626
rect -1287 1438 -1281 1614
rect -1247 1438 -1241 1614
rect -1287 1426 -1241 1438
rect -1129 1614 -1083 1626
rect -1129 1438 -1123 1614
rect -1089 1438 -1083 1614
rect -1129 1426 -1083 1438
rect -971 1614 -925 1626
rect -971 1438 -965 1614
rect -931 1438 -925 1614
rect -971 1426 -925 1438
rect -813 1614 -767 1626
rect -813 1438 -807 1614
rect -773 1438 -767 1614
rect -813 1426 -767 1438
rect -655 1614 -609 1626
rect -655 1438 -649 1614
rect -615 1438 -609 1614
rect -655 1426 -609 1438
rect -497 1614 -451 1626
rect -497 1438 -491 1614
rect -457 1438 -451 1614
rect -497 1426 -451 1438
rect -339 1614 -293 1626
rect -339 1438 -333 1614
rect -299 1438 -293 1614
rect -339 1426 -293 1438
rect -181 1614 -135 1626
rect -181 1438 -175 1614
rect -141 1438 -135 1614
rect -181 1426 -135 1438
rect -23 1614 23 1626
rect -23 1438 -17 1614
rect 17 1438 23 1614
rect -23 1426 23 1438
rect 135 1614 181 1626
rect 135 1438 141 1614
rect 175 1438 181 1614
rect 135 1426 181 1438
rect 293 1614 339 1626
rect 293 1438 299 1614
rect 333 1438 339 1614
rect 293 1426 339 1438
rect 451 1614 497 1626
rect 451 1438 457 1614
rect 491 1438 497 1614
rect 451 1426 497 1438
rect 609 1614 655 1626
rect 609 1438 615 1614
rect 649 1438 655 1614
rect 609 1426 655 1438
rect 767 1614 813 1626
rect 767 1438 773 1614
rect 807 1438 813 1614
rect 767 1426 813 1438
rect 925 1614 971 1626
rect 925 1438 931 1614
rect 965 1438 971 1614
rect 925 1426 971 1438
rect 1083 1614 1129 1626
rect 1083 1438 1089 1614
rect 1123 1438 1129 1614
rect 1083 1426 1129 1438
rect 1241 1614 1287 1626
rect 1241 1438 1247 1614
rect 1281 1438 1287 1614
rect 1241 1426 1287 1438
rect 1399 1614 1445 1626
rect 1399 1438 1405 1614
rect 1439 1438 1445 1614
rect 1399 1426 1445 1438
rect 1557 1614 1603 1626
rect 1557 1438 1563 1614
rect 1597 1438 1603 1614
rect 1557 1426 1603 1438
rect -1547 1379 -1455 1385
rect -1547 1345 -1535 1379
rect -1467 1345 -1455 1379
rect -1547 1339 -1455 1345
rect -1389 1379 -1297 1385
rect -1389 1345 -1377 1379
rect -1309 1345 -1297 1379
rect -1389 1339 -1297 1345
rect -1231 1379 -1139 1385
rect -1231 1345 -1219 1379
rect -1151 1345 -1139 1379
rect -1231 1339 -1139 1345
rect -1073 1379 -981 1385
rect -1073 1345 -1061 1379
rect -993 1345 -981 1379
rect -1073 1339 -981 1345
rect -915 1379 -823 1385
rect -915 1345 -903 1379
rect -835 1345 -823 1379
rect -915 1339 -823 1345
rect -757 1379 -665 1385
rect -757 1345 -745 1379
rect -677 1345 -665 1379
rect -757 1339 -665 1345
rect -599 1379 -507 1385
rect -599 1345 -587 1379
rect -519 1345 -507 1379
rect -599 1339 -507 1345
rect -441 1379 -349 1385
rect -441 1345 -429 1379
rect -361 1345 -349 1379
rect -441 1339 -349 1345
rect -283 1379 -191 1385
rect -283 1345 -271 1379
rect -203 1345 -191 1379
rect -283 1339 -191 1345
rect -125 1379 -33 1385
rect -125 1345 -113 1379
rect -45 1345 -33 1379
rect -125 1339 -33 1345
rect 33 1379 125 1385
rect 33 1345 45 1379
rect 113 1345 125 1379
rect 33 1339 125 1345
rect 191 1379 283 1385
rect 191 1345 203 1379
rect 271 1345 283 1379
rect 191 1339 283 1345
rect 349 1379 441 1385
rect 349 1345 361 1379
rect 429 1345 441 1379
rect 349 1339 441 1345
rect 507 1379 599 1385
rect 507 1345 519 1379
rect 587 1345 599 1379
rect 507 1339 599 1345
rect 665 1379 757 1385
rect 665 1345 677 1379
rect 745 1345 757 1379
rect 665 1339 757 1345
rect 823 1379 915 1385
rect 823 1345 835 1379
rect 903 1345 915 1379
rect 823 1339 915 1345
rect 981 1379 1073 1385
rect 981 1345 993 1379
rect 1061 1345 1073 1379
rect 981 1339 1073 1345
rect 1139 1379 1231 1385
rect 1139 1345 1151 1379
rect 1219 1345 1231 1379
rect 1139 1339 1231 1345
rect 1297 1379 1389 1385
rect 1297 1345 1309 1379
rect 1377 1345 1389 1379
rect 1297 1339 1389 1345
rect 1455 1379 1547 1385
rect 1455 1345 1467 1379
rect 1535 1345 1547 1379
rect 1455 1339 1547 1345
rect -1547 1271 -1455 1277
rect -1547 1237 -1535 1271
rect -1467 1237 -1455 1271
rect -1547 1231 -1455 1237
rect -1389 1271 -1297 1277
rect -1389 1237 -1377 1271
rect -1309 1237 -1297 1271
rect -1389 1231 -1297 1237
rect -1231 1271 -1139 1277
rect -1231 1237 -1219 1271
rect -1151 1237 -1139 1271
rect -1231 1231 -1139 1237
rect -1073 1271 -981 1277
rect -1073 1237 -1061 1271
rect -993 1237 -981 1271
rect -1073 1231 -981 1237
rect -915 1271 -823 1277
rect -915 1237 -903 1271
rect -835 1237 -823 1271
rect -915 1231 -823 1237
rect -757 1271 -665 1277
rect -757 1237 -745 1271
rect -677 1237 -665 1271
rect -757 1231 -665 1237
rect -599 1271 -507 1277
rect -599 1237 -587 1271
rect -519 1237 -507 1271
rect -599 1231 -507 1237
rect -441 1271 -349 1277
rect -441 1237 -429 1271
rect -361 1237 -349 1271
rect -441 1231 -349 1237
rect -283 1271 -191 1277
rect -283 1237 -271 1271
rect -203 1237 -191 1271
rect -283 1231 -191 1237
rect -125 1271 -33 1277
rect -125 1237 -113 1271
rect -45 1237 -33 1271
rect -125 1231 -33 1237
rect 33 1271 125 1277
rect 33 1237 45 1271
rect 113 1237 125 1271
rect 33 1231 125 1237
rect 191 1271 283 1277
rect 191 1237 203 1271
rect 271 1237 283 1271
rect 191 1231 283 1237
rect 349 1271 441 1277
rect 349 1237 361 1271
rect 429 1237 441 1271
rect 349 1231 441 1237
rect 507 1271 599 1277
rect 507 1237 519 1271
rect 587 1237 599 1271
rect 507 1231 599 1237
rect 665 1271 757 1277
rect 665 1237 677 1271
rect 745 1237 757 1271
rect 665 1231 757 1237
rect 823 1271 915 1277
rect 823 1237 835 1271
rect 903 1237 915 1271
rect 823 1231 915 1237
rect 981 1271 1073 1277
rect 981 1237 993 1271
rect 1061 1237 1073 1271
rect 981 1231 1073 1237
rect 1139 1271 1231 1277
rect 1139 1237 1151 1271
rect 1219 1237 1231 1271
rect 1139 1231 1231 1237
rect 1297 1271 1389 1277
rect 1297 1237 1309 1271
rect 1377 1237 1389 1271
rect 1297 1231 1389 1237
rect 1455 1271 1547 1277
rect 1455 1237 1467 1271
rect 1535 1237 1547 1271
rect 1455 1231 1547 1237
rect -1603 1178 -1557 1190
rect -1603 1002 -1597 1178
rect -1563 1002 -1557 1178
rect -1603 990 -1557 1002
rect -1445 1178 -1399 1190
rect -1445 1002 -1439 1178
rect -1405 1002 -1399 1178
rect -1445 990 -1399 1002
rect -1287 1178 -1241 1190
rect -1287 1002 -1281 1178
rect -1247 1002 -1241 1178
rect -1287 990 -1241 1002
rect -1129 1178 -1083 1190
rect -1129 1002 -1123 1178
rect -1089 1002 -1083 1178
rect -1129 990 -1083 1002
rect -971 1178 -925 1190
rect -971 1002 -965 1178
rect -931 1002 -925 1178
rect -971 990 -925 1002
rect -813 1178 -767 1190
rect -813 1002 -807 1178
rect -773 1002 -767 1178
rect -813 990 -767 1002
rect -655 1178 -609 1190
rect -655 1002 -649 1178
rect -615 1002 -609 1178
rect -655 990 -609 1002
rect -497 1178 -451 1190
rect -497 1002 -491 1178
rect -457 1002 -451 1178
rect -497 990 -451 1002
rect -339 1178 -293 1190
rect -339 1002 -333 1178
rect -299 1002 -293 1178
rect -339 990 -293 1002
rect -181 1178 -135 1190
rect -181 1002 -175 1178
rect -141 1002 -135 1178
rect -181 990 -135 1002
rect -23 1178 23 1190
rect -23 1002 -17 1178
rect 17 1002 23 1178
rect -23 990 23 1002
rect 135 1178 181 1190
rect 135 1002 141 1178
rect 175 1002 181 1178
rect 135 990 181 1002
rect 293 1178 339 1190
rect 293 1002 299 1178
rect 333 1002 339 1178
rect 293 990 339 1002
rect 451 1178 497 1190
rect 451 1002 457 1178
rect 491 1002 497 1178
rect 451 990 497 1002
rect 609 1178 655 1190
rect 609 1002 615 1178
rect 649 1002 655 1178
rect 609 990 655 1002
rect 767 1178 813 1190
rect 767 1002 773 1178
rect 807 1002 813 1178
rect 767 990 813 1002
rect 925 1178 971 1190
rect 925 1002 931 1178
rect 965 1002 971 1178
rect 925 990 971 1002
rect 1083 1178 1129 1190
rect 1083 1002 1089 1178
rect 1123 1002 1129 1178
rect 1083 990 1129 1002
rect 1241 1178 1287 1190
rect 1241 1002 1247 1178
rect 1281 1002 1287 1178
rect 1241 990 1287 1002
rect 1399 1178 1445 1190
rect 1399 1002 1405 1178
rect 1439 1002 1445 1178
rect 1399 990 1445 1002
rect 1557 1178 1603 1190
rect 1557 1002 1563 1178
rect 1597 1002 1603 1178
rect 1557 990 1603 1002
rect -1547 943 -1455 949
rect -1547 909 -1535 943
rect -1467 909 -1455 943
rect -1547 903 -1455 909
rect -1389 943 -1297 949
rect -1389 909 -1377 943
rect -1309 909 -1297 943
rect -1389 903 -1297 909
rect -1231 943 -1139 949
rect -1231 909 -1219 943
rect -1151 909 -1139 943
rect -1231 903 -1139 909
rect -1073 943 -981 949
rect -1073 909 -1061 943
rect -993 909 -981 943
rect -1073 903 -981 909
rect -915 943 -823 949
rect -915 909 -903 943
rect -835 909 -823 943
rect -915 903 -823 909
rect -757 943 -665 949
rect -757 909 -745 943
rect -677 909 -665 943
rect -757 903 -665 909
rect -599 943 -507 949
rect -599 909 -587 943
rect -519 909 -507 943
rect -599 903 -507 909
rect -441 943 -349 949
rect -441 909 -429 943
rect -361 909 -349 943
rect -441 903 -349 909
rect -283 943 -191 949
rect -283 909 -271 943
rect -203 909 -191 943
rect -283 903 -191 909
rect -125 943 -33 949
rect -125 909 -113 943
rect -45 909 -33 943
rect -125 903 -33 909
rect 33 943 125 949
rect 33 909 45 943
rect 113 909 125 943
rect 33 903 125 909
rect 191 943 283 949
rect 191 909 203 943
rect 271 909 283 943
rect 191 903 283 909
rect 349 943 441 949
rect 349 909 361 943
rect 429 909 441 943
rect 349 903 441 909
rect 507 943 599 949
rect 507 909 519 943
rect 587 909 599 943
rect 507 903 599 909
rect 665 943 757 949
rect 665 909 677 943
rect 745 909 757 943
rect 665 903 757 909
rect 823 943 915 949
rect 823 909 835 943
rect 903 909 915 943
rect 823 903 915 909
rect 981 943 1073 949
rect 981 909 993 943
rect 1061 909 1073 943
rect 981 903 1073 909
rect 1139 943 1231 949
rect 1139 909 1151 943
rect 1219 909 1231 943
rect 1139 903 1231 909
rect 1297 943 1389 949
rect 1297 909 1309 943
rect 1377 909 1389 943
rect 1297 903 1389 909
rect 1455 943 1547 949
rect 1455 909 1467 943
rect 1535 909 1547 943
rect 1455 903 1547 909
rect -1547 835 -1455 841
rect -1547 801 -1535 835
rect -1467 801 -1455 835
rect -1547 795 -1455 801
rect -1389 835 -1297 841
rect -1389 801 -1377 835
rect -1309 801 -1297 835
rect -1389 795 -1297 801
rect -1231 835 -1139 841
rect -1231 801 -1219 835
rect -1151 801 -1139 835
rect -1231 795 -1139 801
rect -1073 835 -981 841
rect -1073 801 -1061 835
rect -993 801 -981 835
rect -1073 795 -981 801
rect -915 835 -823 841
rect -915 801 -903 835
rect -835 801 -823 835
rect -915 795 -823 801
rect -757 835 -665 841
rect -757 801 -745 835
rect -677 801 -665 835
rect -757 795 -665 801
rect -599 835 -507 841
rect -599 801 -587 835
rect -519 801 -507 835
rect -599 795 -507 801
rect -441 835 -349 841
rect -441 801 -429 835
rect -361 801 -349 835
rect -441 795 -349 801
rect -283 835 -191 841
rect -283 801 -271 835
rect -203 801 -191 835
rect -283 795 -191 801
rect -125 835 -33 841
rect -125 801 -113 835
rect -45 801 -33 835
rect -125 795 -33 801
rect 33 835 125 841
rect 33 801 45 835
rect 113 801 125 835
rect 33 795 125 801
rect 191 835 283 841
rect 191 801 203 835
rect 271 801 283 835
rect 191 795 283 801
rect 349 835 441 841
rect 349 801 361 835
rect 429 801 441 835
rect 349 795 441 801
rect 507 835 599 841
rect 507 801 519 835
rect 587 801 599 835
rect 507 795 599 801
rect 665 835 757 841
rect 665 801 677 835
rect 745 801 757 835
rect 665 795 757 801
rect 823 835 915 841
rect 823 801 835 835
rect 903 801 915 835
rect 823 795 915 801
rect 981 835 1073 841
rect 981 801 993 835
rect 1061 801 1073 835
rect 981 795 1073 801
rect 1139 835 1231 841
rect 1139 801 1151 835
rect 1219 801 1231 835
rect 1139 795 1231 801
rect 1297 835 1389 841
rect 1297 801 1309 835
rect 1377 801 1389 835
rect 1297 795 1389 801
rect 1455 835 1547 841
rect 1455 801 1467 835
rect 1535 801 1547 835
rect 1455 795 1547 801
rect -1603 742 -1557 754
rect -1603 566 -1597 742
rect -1563 566 -1557 742
rect -1603 554 -1557 566
rect -1445 742 -1399 754
rect -1445 566 -1439 742
rect -1405 566 -1399 742
rect -1445 554 -1399 566
rect -1287 742 -1241 754
rect -1287 566 -1281 742
rect -1247 566 -1241 742
rect -1287 554 -1241 566
rect -1129 742 -1083 754
rect -1129 566 -1123 742
rect -1089 566 -1083 742
rect -1129 554 -1083 566
rect -971 742 -925 754
rect -971 566 -965 742
rect -931 566 -925 742
rect -971 554 -925 566
rect -813 742 -767 754
rect -813 566 -807 742
rect -773 566 -767 742
rect -813 554 -767 566
rect -655 742 -609 754
rect -655 566 -649 742
rect -615 566 -609 742
rect -655 554 -609 566
rect -497 742 -451 754
rect -497 566 -491 742
rect -457 566 -451 742
rect -497 554 -451 566
rect -339 742 -293 754
rect -339 566 -333 742
rect -299 566 -293 742
rect -339 554 -293 566
rect -181 742 -135 754
rect -181 566 -175 742
rect -141 566 -135 742
rect -181 554 -135 566
rect -23 742 23 754
rect -23 566 -17 742
rect 17 566 23 742
rect -23 554 23 566
rect 135 742 181 754
rect 135 566 141 742
rect 175 566 181 742
rect 135 554 181 566
rect 293 742 339 754
rect 293 566 299 742
rect 333 566 339 742
rect 293 554 339 566
rect 451 742 497 754
rect 451 566 457 742
rect 491 566 497 742
rect 451 554 497 566
rect 609 742 655 754
rect 609 566 615 742
rect 649 566 655 742
rect 609 554 655 566
rect 767 742 813 754
rect 767 566 773 742
rect 807 566 813 742
rect 767 554 813 566
rect 925 742 971 754
rect 925 566 931 742
rect 965 566 971 742
rect 925 554 971 566
rect 1083 742 1129 754
rect 1083 566 1089 742
rect 1123 566 1129 742
rect 1083 554 1129 566
rect 1241 742 1287 754
rect 1241 566 1247 742
rect 1281 566 1287 742
rect 1241 554 1287 566
rect 1399 742 1445 754
rect 1399 566 1405 742
rect 1439 566 1445 742
rect 1399 554 1445 566
rect 1557 742 1603 754
rect 1557 566 1563 742
rect 1597 566 1603 742
rect 1557 554 1603 566
rect -1547 507 -1455 513
rect -1547 473 -1535 507
rect -1467 473 -1455 507
rect -1547 467 -1455 473
rect -1389 507 -1297 513
rect -1389 473 -1377 507
rect -1309 473 -1297 507
rect -1389 467 -1297 473
rect -1231 507 -1139 513
rect -1231 473 -1219 507
rect -1151 473 -1139 507
rect -1231 467 -1139 473
rect -1073 507 -981 513
rect -1073 473 -1061 507
rect -993 473 -981 507
rect -1073 467 -981 473
rect -915 507 -823 513
rect -915 473 -903 507
rect -835 473 -823 507
rect -915 467 -823 473
rect -757 507 -665 513
rect -757 473 -745 507
rect -677 473 -665 507
rect -757 467 -665 473
rect -599 507 -507 513
rect -599 473 -587 507
rect -519 473 -507 507
rect -599 467 -507 473
rect -441 507 -349 513
rect -441 473 -429 507
rect -361 473 -349 507
rect -441 467 -349 473
rect -283 507 -191 513
rect -283 473 -271 507
rect -203 473 -191 507
rect -283 467 -191 473
rect -125 507 -33 513
rect -125 473 -113 507
rect -45 473 -33 507
rect -125 467 -33 473
rect 33 507 125 513
rect 33 473 45 507
rect 113 473 125 507
rect 33 467 125 473
rect 191 507 283 513
rect 191 473 203 507
rect 271 473 283 507
rect 191 467 283 473
rect 349 507 441 513
rect 349 473 361 507
rect 429 473 441 507
rect 349 467 441 473
rect 507 507 599 513
rect 507 473 519 507
rect 587 473 599 507
rect 507 467 599 473
rect 665 507 757 513
rect 665 473 677 507
rect 745 473 757 507
rect 665 467 757 473
rect 823 507 915 513
rect 823 473 835 507
rect 903 473 915 507
rect 823 467 915 473
rect 981 507 1073 513
rect 981 473 993 507
rect 1061 473 1073 507
rect 981 467 1073 473
rect 1139 507 1231 513
rect 1139 473 1151 507
rect 1219 473 1231 507
rect 1139 467 1231 473
rect 1297 507 1389 513
rect 1297 473 1309 507
rect 1377 473 1389 507
rect 1297 467 1389 473
rect 1455 507 1547 513
rect 1455 473 1467 507
rect 1535 473 1547 507
rect 1455 467 1547 473
rect -1547 399 -1455 405
rect -1547 365 -1535 399
rect -1467 365 -1455 399
rect -1547 359 -1455 365
rect -1389 399 -1297 405
rect -1389 365 -1377 399
rect -1309 365 -1297 399
rect -1389 359 -1297 365
rect -1231 399 -1139 405
rect -1231 365 -1219 399
rect -1151 365 -1139 399
rect -1231 359 -1139 365
rect -1073 399 -981 405
rect -1073 365 -1061 399
rect -993 365 -981 399
rect -1073 359 -981 365
rect -915 399 -823 405
rect -915 365 -903 399
rect -835 365 -823 399
rect -915 359 -823 365
rect -757 399 -665 405
rect -757 365 -745 399
rect -677 365 -665 399
rect -757 359 -665 365
rect -599 399 -507 405
rect -599 365 -587 399
rect -519 365 -507 399
rect -599 359 -507 365
rect -441 399 -349 405
rect -441 365 -429 399
rect -361 365 -349 399
rect -441 359 -349 365
rect -283 399 -191 405
rect -283 365 -271 399
rect -203 365 -191 399
rect -283 359 -191 365
rect -125 399 -33 405
rect -125 365 -113 399
rect -45 365 -33 399
rect -125 359 -33 365
rect 33 399 125 405
rect 33 365 45 399
rect 113 365 125 399
rect 33 359 125 365
rect 191 399 283 405
rect 191 365 203 399
rect 271 365 283 399
rect 191 359 283 365
rect 349 399 441 405
rect 349 365 361 399
rect 429 365 441 399
rect 349 359 441 365
rect 507 399 599 405
rect 507 365 519 399
rect 587 365 599 399
rect 507 359 599 365
rect 665 399 757 405
rect 665 365 677 399
rect 745 365 757 399
rect 665 359 757 365
rect 823 399 915 405
rect 823 365 835 399
rect 903 365 915 399
rect 823 359 915 365
rect 981 399 1073 405
rect 981 365 993 399
rect 1061 365 1073 399
rect 981 359 1073 365
rect 1139 399 1231 405
rect 1139 365 1151 399
rect 1219 365 1231 399
rect 1139 359 1231 365
rect 1297 399 1389 405
rect 1297 365 1309 399
rect 1377 365 1389 399
rect 1297 359 1389 365
rect 1455 399 1547 405
rect 1455 365 1467 399
rect 1535 365 1547 399
rect 1455 359 1547 365
rect -1603 306 -1557 318
rect -1603 130 -1597 306
rect -1563 130 -1557 306
rect -1603 118 -1557 130
rect -1445 306 -1399 318
rect -1445 130 -1439 306
rect -1405 130 -1399 306
rect -1445 118 -1399 130
rect -1287 306 -1241 318
rect -1287 130 -1281 306
rect -1247 130 -1241 306
rect -1287 118 -1241 130
rect -1129 306 -1083 318
rect -1129 130 -1123 306
rect -1089 130 -1083 306
rect -1129 118 -1083 130
rect -971 306 -925 318
rect -971 130 -965 306
rect -931 130 -925 306
rect -971 118 -925 130
rect -813 306 -767 318
rect -813 130 -807 306
rect -773 130 -767 306
rect -813 118 -767 130
rect -655 306 -609 318
rect -655 130 -649 306
rect -615 130 -609 306
rect -655 118 -609 130
rect -497 306 -451 318
rect -497 130 -491 306
rect -457 130 -451 306
rect -497 118 -451 130
rect -339 306 -293 318
rect -339 130 -333 306
rect -299 130 -293 306
rect -339 118 -293 130
rect -181 306 -135 318
rect -181 130 -175 306
rect -141 130 -135 306
rect -181 118 -135 130
rect -23 306 23 318
rect -23 130 -17 306
rect 17 130 23 306
rect -23 118 23 130
rect 135 306 181 318
rect 135 130 141 306
rect 175 130 181 306
rect 135 118 181 130
rect 293 306 339 318
rect 293 130 299 306
rect 333 130 339 306
rect 293 118 339 130
rect 451 306 497 318
rect 451 130 457 306
rect 491 130 497 306
rect 451 118 497 130
rect 609 306 655 318
rect 609 130 615 306
rect 649 130 655 306
rect 609 118 655 130
rect 767 306 813 318
rect 767 130 773 306
rect 807 130 813 306
rect 767 118 813 130
rect 925 306 971 318
rect 925 130 931 306
rect 965 130 971 306
rect 925 118 971 130
rect 1083 306 1129 318
rect 1083 130 1089 306
rect 1123 130 1129 306
rect 1083 118 1129 130
rect 1241 306 1287 318
rect 1241 130 1247 306
rect 1281 130 1287 306
rect 1241 118 1287 130
rect 1399 306 1445 318
rect 1399 130 1405 306
rect 1439 130 1445 306
rect 1399 118 1445 130
rect 1557 306 1603 318
rect 1557 130 1563 306
rect 1597 130 1603 306
rect 1557 118 1603 130
rect -1547 71 -1455 77
rect -1547 37 -1535 71
rect -1467 37 -1455 71
rect -1547 31 -1455 37
rect -1389 71 -1297 77
rect -1389 37 -1377 71
rect -1309 37 -1297 71
rect -1389 31 -1297 37
rect -1231 71 -1139 77
rect -1231 37 -1219 71
rect -1151 37 -1139 71
rect -1231 31 -1139 37
rect -1073 71 -981 77
rect -1073 37 -1061 71
rect -993 37 -981 71
rect -1073 31 -981 37
rect -915 71 -823 77
rect -915 37 -903 71
rect -835 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 835 71
rect 903 37 915 71
rect 823 31 915 37
rect 981 71 1073 77
rect 981 37 993 71
rect 1061 37 1073 71
rect 981 31 1073 37
rect 1139 71 1231 77
rect 1139 37 1151 71
rect 1219 37 1231 71
rect 1139 31 1231 37
rect 1297 71 1389 77
rect 1297 37 1309 71
rect 1377 37 1389 71
rect 1297 31 1389 37
rect 1455 71 1547 77
rect 1455 37 1467 71
rect 1535 37 1547 71
rect 1455 31 1547 37
rect -1547 -37 -1455 -31
rect -1547 -71 -1535 -37
rect -1467 -71 -1455 -37
rect -1547 -77 -1455 -71
rect -1389 -37 -1297 -31
rect -1389 -71 -1377 -37
rect -1309 -71 -1297 -37
rect -1389 -77 -1297 -71
rect -1231 -37 -1139 -31
rect -1231 -71 -1219 -37
rect -1151 -71 -1139 -37
rect -1231 -77 -1139 -71
rect -1073 -37 -981 -31
rect -1073 -71 -1061 -37
rect -993 -71 -981 -37
rect -1073 -77 -981 -71
rect -915 -37 -823 -31
rect -915 -71 -903 -37
rect -835 -71 -823 -37
rect -915 -77 -823 -71
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect 823 -37 915 -31
rect 823 -71 835 -37
rect 903 -71 915 -37
rect 823 -77 915 -71
rect 981 -37 1073 -31
rect 981 -71 993 -37
rect 1061 -71 1073 -37
rect 981 -77 1073 -71
rect 1139 -37 1231 -31
rect 1139 -71 1151 -37
rect 1219 -71 1231 -37
rect 1139 -77 1231 -71
rect 1297 -37 1389 -31
rect 1297 -71 1309 -37
rect 1377 -71 1389 -37
rect 1297 -77 1389 -71
rect 1455 -37 1547 -31
rect 1455 -71 1467 -37
rect 1535 -71 1547 -37
rect 1455 -77 1547 -71
rect -1603 -130 -1557 -118
rect -1603 -306 -1597 -130
rect -1563 -306 -1557 -130
rect -1603 -318 -1557 -306
rect -1445 -130 -1399 -118
rect -1445 -306 -1439 -130
rect -1405 -306 -1399 -130
rect -1445 -318 -1399 -306
rect -1287 -130 -1241 -118
rect -1287 -306 -1281 -130
rect -1247 -306 -1241 -130
rect -1287 -318 -1241 -306
rect -1129 -130 -1083 -118
rect -1129 -306 -1123 -130
rect -1089 -306 -1083 -130
rect -1129 -318 -1083 -306
rect -971 -130 -925 -118
rect -971 -306 -965 -130
rect -931 -306 -925 -130
rect -971 -318 -925 -306
rect -813 -130 -767 -118
rect -813 -306 -807 -130
rect -773 -306 -767 -130
rect -813 -318 -767 -306
rect -655 -130 -609 -118
rect -655 -306 -649 -130
rect -615 -306 -609 -130
rect -655 -318 -609 -306
rect -497 -130 -451 -118
rect -497 -306 -491 -130
rect -457 -306 -451 -130
rect -497 -318 -451 -306
rect -339 -130 -293 -118
rect -339 -306 -333 -130
rect -299 -306 -293 -130
rect -339 -318 -293 -306
rect -181 -130 -135 -118
rect -181 -306 -175 -130
rect -141 -306 -135 -130
rect -181 -318 -135 -306
rect -23 -130 23 -118
rect -23 -306 -17 -130
rect 17 -306 23 -130
rect -23 -318 23 -306
rect 135 -130 181 -118
rect 135 -306 141 -130
rect 175 -306 181 -130
rect 135 -318 181 -306
rect 293 -130 339 -118
rect 293 -306 299 -130
rect 333 -306 339 -130
rect 293 -318 339 -306
rect 451 -130 497 -118
rect 451 -306 457 -130
rect 491 -306 497 -130
rect 451 -318 497 -306
rect 609 -130 655 -118
rect 609 -306 615 -130
rect 649 -306 655 -130
rect 609 -318 655 -306
rect 767 -130 813 -118
rect 767 -306 773 -130
rect 807 -306 813 -130
rect 767 -318 813 -306
rect 925 -130 971 -118
rect 925 -306 931 -130
rect 965 -306 971 -130
rect 925 -318 971 -306
rect 1083 -130 1129 -118
rect 1083 -306 1089 -130
rect 1123 -306 1129 -130
rect 1083 -318 1129 -306
rect 1241 -130 1287 -118
rect 1241 -306 1247 -130
rect 1281 -306 1287 -130
rect 1241 -318 1287 -306
rect 1399 -130 1445 -118
rect 1399 -306 1405 -130
rect 1439 -306 1445 -130
rect 1399 -318 1445 -306
rect 1557 -130 1603 -118
rect 1557 -306 1563 -130
rect 1597 -306 1603 -130
rect 1557 -318 1603 -306
rect -1547 -365 -1455 -359
rect -1547 -399 -1535 -365
rect -1467 -399 -1455 -365
rect -1547 -405 -1455 -399
rect -1389 -365 -1297 -359
rect -1389 -399 -1377 -365
rect -1309 -399 -1297 -365
rect -1389 -405 -1297 -399
rect -1231 -365 -1139 -359
rect -1231 -399 -1219 -365
rect -1151 -399 -1139 -365
rect -1231 -405 -1139 -399
rect -1073 -365 -981 -359
rect -1073 -399 -1061 -365
rect -993 -399 -981 -365
rect -1073 -405 -981 -399
rect -915 -365 -823 -359
rect -915 -399 -903 -365
rect -835 -399 -823 -365
rect -915 -405 -823 -399
rect -757 -365 -665 -359
rect -757 -399 -745 -365
rect -677 -399 -665 -365
rect -757 -405 -665 -399
rect -599 -365 -507 -359
rect -599 -399 -587 -365
rect -519 -399 -507 -365
rect -599 -405 -507 -399
rect -441 -365 -349 -359
rect -441 -399 -429 -365
rect -361 -399 -349 -365
rect -441 -405 -349 -399
rect -283 -365 -191 -359
rect -283 -399 -271 -365
rect -203 -399 -191 -365
rect -283 -405 -191 -399
rect -125 -365 -33 -359
rect -125 -399 -113 -365
rect -45 -399 -33 -365
rect -125 -405 -33 -399
rect 33 -365 125 -359
rect 33 -399 45 -365
rect 113 -399 125 -365
rect 33 -405 125 -399
rect 191 -365 283 -359
rect 191 -399 203 -365
rect 271 -399 283 -365
rect 191 -405 283 -399
rect 349 -365 441 -359
rect 349 -399 361 -365
rect 429 -399 441 -365
rect 349 -405 441 -399
rect 507 -365 599 -359
rect 507 -399 519 -365
rect 587 -399 599 -365
rect 507 -405 599 -399
rect 665 -365 757 -359
rect 665 -399 677 -365
rect 745 -399 757 -365
rect 665 -405 757 -399
rect 823 -365 915 -359
rect 823 -399 835 -365
rect 903 -399 915 -365
rect 823 -405 915 -399
rect 981 -365 1073 -359
rect 981 -399 993 -365
rect 1061 -399 1073 -365
rect 981 -405 1073 -399
rect 1139 -365 1231 -359
rect 1139 -399 1151 -365
rect 1219 -399 1231 -365
rect 1139 -405 1231 -399
rect 1297 -365 1389 -359
rect 1297 -399 1309 -365
rect 1377 -399 1389 -365
rect 1297 -405 1389 -399
rect 1455 -365 1547 -359
rect 1455 -399 1467 -365
rect 1535 -399 1547 -365
rect 1455 -405 1547 -399
rect -1547 -473 -1455 -467
rect -1547 -507 -1535 -473
rect -1467 -507 -1455 -473
rect -1547 -513 -1455 -507
rect -1389 -473 -1297 -467
rect -1389 -507 -1377 -473
rect -1309 -507 -1297 -473
rect -1389 -513 -1297 -507
rect -1231 -473 -1139 -467
rect -1231 -507 -1219 -473
rect -1151 -507 -1139 -473
rect -1231 -513 -1139 -507
rect -1073 -473 -981 -467
rect -1073 -507 -1061 -473
rect -993 -507 -981 -473
rect -1073 -513 -981 -507
rect -915 -473 -823 -467
rect -915 -507 -903 -473
rect -835 -507 -823 -473
rect -915 -513 -823 -507
rect -757 -473 -665 -467
rect -757 -507 -745 -473
rect -677 -507 -665 -473
rect -757 -513 -665 -507
rect -599 -473 -507 -467
rect -599 -507 -587 -473
rect -519 -507 -507 -473
rect -599 -513 -507 -507
rect -441 -473 -349 -467
rect -441 -507 -429 -473
rect -361 -507 -349 -473
rect -441 -513 -349 -507
rect -283 -473 -191 -467
rect -283 -507 -271 -473
rect -203 -507 -191 -473
rect -283 -513 -191 -507
rect -125 -473 -33 -467
rect -125 -507 -113 -473
rect -45 -507 -33 -473
rect -125 -513 -33 -507
rect 33 -473 125 -467
rect 33 -507 45 -473
rect 113 -507 125 -473
rect 33 -513 125 -507
rect 191 -473 283 -467
rect 191 -507 203 -473
rect 271 -507 283 -473
rect 191 -513 283 -507
rect 349 -473 441 -467
rect 349 -507 361 -473
rect 429 -507 441 -473
rect 349 -513 441 -507
rect 507 -473 599 -467
rect 507 -507 519 -473
rect 587 -507 599 -473
rect 507 -513 599 -507
rect 665 -473 757 -467
rect 665 -507 677 -473
rect 745 -507 757 -473
rect 665 -513 757 -507
rect 823 -473 915 -467
rect 823 -507 835 -473
rect 903 -507 915 -473
rect 823 -513 915 -507
rect 981 -473 1073 -467
rect 981 -507 993 -473
rect 1061 -507 1073 -473
rect 981 -513 1073 -507
rect 1139 -473 1231 -467
rect 1139 -507 1151 -473
rect 1219 -507 1231 -473
rect 1139 -513 1231 -507
rect 1297 -473 1389 -467
rect 1297 -507 1309 -473
rect 1377 -507 1389 -473
rect 1297 -513 1389 -507
rect 1455 -473 1547 -467
rect 1455 -507 1467 -473
rect 1535 -507 1547 -473
rect 1455 -513 1547 -507
rect -1603 -566 -1557 -554
rect -1603 -742 -1597 -566
rect -1563 -742 -1557 -566
rect -1603 -754 -1557 -742
rect -1445 -566 -1399 -554
rect -1445 -742 -1439 -566
rect -1405 -742 -1399 -566
rect -1445 -754 -1399 -742
rect -1287 -566 -1241 -554
rect -1287 -742 -1281 -566
rect -1247 -742 -1241 -566
rect -1287 -754 -1241 -742
rect -1129 -566 -1083 -554
rect -1129 -742 -1123 -566
rect -1089 -742 -1083 -566
rect -1129 -754 -1083 -742
rect -971 -566 -925 -554
rect -971 -742 -965 -566
rect -931 -742 -925 -566
rect -971 -754 -925 -742
rect -813 -566 -767 -554
rect -813 -742 -807 -566
rect -773 -742 -767 -566
rect -813 -754 -767 -742
rect -655 -566 -609 -554
rect -655 -742 -649 -566
rect -615 -742 -609 -566
rect -655 -754 -609 -742
rect -497 -566 -451 -554
rect -497 -742 -491 -566
rect -457 -742 -451 -566
rect -497 -754 -451 -742
rect -339 -566 -293 -554
rect -339 -742 -333 -566
rect -299 -742 -293 -566
rect -339 -754 -293 -742
rect -181 -566 -135 -554
rect -181 -742 -175 -566
rect -141 -742 -135 -566
rect -181 -754 -135 -742
rect -23 -566 23 -554
rect -23 -742 -17 -566
rect 17 -742 23 -566
rect -23 -754 23 -742
rect 135 -566 181 -554
rect 135 -742 141 -566
rect 175 -742 181 -566
rect 135 -754 181 -742
rect 293 -566 339 -554
rect 293 -742 299 -566
rect 333 -742 339 -566
rect 293 -754 339 -742
rect 451 -566 497 -554
rect 451 -742 457 -566
rect 491 -742 497 -566
rect 451 -754 497 -742
rect 609 -566 655 -554
rect 609 -742 615 -566
rect 649 -742 655 -566
rect 609 -754 655 -742
rect 767 -566 813 -554
rect 767 -742 773 -566
rect 807 -742 813 -566
rect 767 -754 813 -742
rect 925 -566 971 -554
rect 925 -742 931 -566
rect 965 -742 971 -566
rect 925 -754 971 -742
rect 1083 -566 1129 -554
rect 1083 -742 1089 -566
rect 1123 -742 1129 -566
rect 1083 -754 1129 -742
rect 1241 -566 1287 -554
rect 1241 -742 1247 -566
rect 1281 -742 1287 -566
rect 1241 -754 1287 -742
rect 1399 -566 1445 -554
rect 1399 -742 1405 -566
rect 1439 -742 1445 -566
rect 1399 -754 1445 -742
rect 1557 -566 1603 -554
rect 1557 -742 1563 -566
rect 1597 -742 1603 -566
rect 1557 -754 1603 -742
rect -1547 -801 -1455 -795
rect -1547 -835 -1535 -801
rect -1467 -835 -1455 -801
rect -1547 -841 -1455 -835
rect -1389 -801 -1297 -795
rect -1389 -835 -1377 -801
rect -1309 -835 -1297 -801
rect -1389 -841 -1297 -835
rect -1231 -801 -1139 -795
rect -1231 -835 -1219 -801
rect -1151 -835 -1139 -801
rect -1231 -841 -1139 -835
rect -1073 -801 -981 -795
rect -1073 -835 -1061 -801
rect -993 -835 -981 -801
rect -1073 -841 -981 -835
rect -915 -801 -823 -795
rect -915 -835 -903 -801
rect -835 -835 -823 -801
rect -915 -841 -823 -835
rect -757 -801 -665 -795
rect -757 -835 -745 -801
rect -677 -835 -665 -801
rect -757 -841 -665 -835
rect -599 -801 -507 -795
rect -599 -835 -587 -801
rect -519 -835 -507 -801
rect -599 -841 -507 -835
rect -441 -801 -349 -795
rect -441 -835 -429 -801
rect -361 -835 -349 -801
rect -441 -841 -349 -835
rect -283 -801 -191 -795
rect -283 -835 -271 -801
rect -203 -835 -191 -801
rect -283 -841 -191 -835
rect -125 -801 -33 -795
rect -125 -835 -113 -801
rect -45 -835 -33 -801
rect -125 -841 -33 -835
rect 33 -801 125 -795
rect 33 -835 45 -801
rect 113 -835 125 -801
rect 33 -841 125 -835
rect 191 -801 283 -795
rect 191 -835 203 -801
rect 271 -835 283 -801
rect 191 -841 283 -835
rect 349 -801 441 -795
rect 349 -835 361 -801
rect 429 -835 441 -801
rect 349 -841 441 -835
rect 507 -801 599 -795
rect 507 -835 519 -801
rect 587 -835 599 -801
rect 507 -841 599 -835
rect 665 -801 757 -795
rect 665 -835 677 -801
rect 745 -835 757 -801
rect 665 -841 757 -835
rect 823 -801 915 -795
rect 823 -835 835 -801
rect 903 -835 915 -801
rect 823 -841 915 -835
rect 981 -801 1073 -795
rect 981 -835 993 -801
rect 1061 -835 1073 -801
rect 981 -841 1073 -835
rect 1139 -801 1231 -795
rect 1139 -835 1151 -801
rect 1219 -835 1231 -801
rect 1139 -841 1231 -835
rect 1297 -801 1389 -795
rect 1297 -835 1309 -801
rect 1377 -835 1389 -801
rect 1297 -841 1389 -835
rect 1455 -801 1547 -795
rect 1455 -835 1467 -801
rect 1535 -835 1547 -801
rect 1455 -841 1547 -835
rect -1547 -909 -1455 -903
rect -1547 -943 -1535 -909
rect -1467 -943 -1455 -909
rect -1547 -949 -1455 -943
rect -1389 -909 -1297 -903
rect -1389 -943 -1377 -909
rect -1309 -943 -1297 -909
rect -1389 -949 -1297 -943
rect -1231 -909 -1139 -903
rect -1231 -943 -1219 -909
rect -1151 -943 -1139 -909
rect -1231 -949 -1139 -943
rect -1073 -909 -981 -903
rect -1073 -943 -1061 -909
rect -993 -943 -981 -909
rect -1073 -949 -981 -943
rect -915 -909 -823 -903
rect -915 -943 -903 -909
rect -835 -943 -823 -909
rect -915 -949 -823 -943
rect -757 -909 -665 -903
rect -757 -943 -745 -909
rect -677 -943 -665 -909
rect -757 -949 -665 -943
rect -599 -909 -507 -903
rect -599 -943 -587 -909
rect -519 -943 -507 -909
rect -599 -949 -507 -943
rect -441 -909 -349 -903
rect -441 -943 -429 -909
rect -361 -943 -349 -909
rect -441 -949 -349 -943
rect -283 -909 -191 -903
rect -283 -943 -271 -909
rect -203 -943 -191 -909
rect -283 -949 -191 -943
rect -125 -909 -33 -903
rect -125 -943 -113 -909
rect -45 -943 -33 -909
rect -125 -949 -33 -943
rect 33 -909 125 -903
rect 33 -943 45 -909
rect 113 -943 125 -909
rect 33 -949 125 -943
rect 191 -909 283 -903
rect 191 -943 203 -909
rect 271 -943 283 -909
rect 191 -949 283 -943
rect 349 -909 441 -903
rect 349 -943 361 -909
rect 429 -943 441 -909
rect 349 -949 441 -943
rect 507 -909 599 -903
rect 507 -943 519 -909
rect 587 -943 599 -909
rect 507 -949 599 -943
rect 665 -909 757 -903
rect 665 -943 677 -909
rect 745 -943 757 -909
rect 665 -949 757 -943
rect 823 -909 915 -903
rect 823 -943 835 -909
rect 903 -943 915 -909
rect 823 -949 915 -943
rect 981 -909 1073 -903
rect 981 -943 993 -909
rect 1061 -943 1073 -909
rect 981 -949 1073 -943
rect 1139 -909 1231 -903
rect 1139 -943 1151 -909
rect 1219 -943 1231 -909
rect 1139 -949 1231 -943
rect 1297 -909 1389 -903
rect 1297 -943 1309 -909
rect 1377 -943 1389 -909
rect 1297 -949 1389 -943
rect 1455 -909 1547 -903
rect 1455 -943 1467 -909
rect 1535 -943 1547 -909
rect 1455 -949 1547 -943
rect -1603 -1002 -1557 -990
rect -1603 -1178 -1597 -1002
rect -1563 -1178 -1557 -1002
rect -1603 -1190 -1557 -1178
rect -1445 -1002 -1399 -990
rect -1445 -1178 -1439 -1002
rect -1405 -1178 -1399 -1002
rect -1445 -1190 -1399 -1178
rect -1287 -1002 -1241 -990
rect -1287 -1178 -1281 -1002
rect -1247 -1178 -1241 -1002
rect -1287 -1190 -1241 -1178
rect -1129 -1002 -1083 -990
rect -1129 -1178 -1123 -1002
rect -1089 -1178 -1083 -1002
rect -1129 -1190 -1083 -1178
rect -971 -1002 -925 -990
rect -971 -1178 -965 -1002
rect -931 -1178 -925 -1002
rect -971 -1190 -925 -1178
rect -813 -1002 -767 -990
rect -813 -1178 -807 -1002
rect -773 -1178 -767 -1002
rect -813 -1190 -767 -1178
rect -655 -1002 -609 -990
rect -655 -1178 -649 -1002
rect -615 -1178 -609 -1002
rect -655 -1190 -609 -1178
rect -497 -1002 -451 -990
rect -497 -1178 -491 -1002
rect -457 -1178 -451 -1002
rect -497 -1190 -451 -1178
rect -339 -1002 -293 -990
rect -339 -1178 -333 -1002
rect -299 -1178 -293 -1002
rect -339 -1190 -293 -1178
rect -181 -1002 -135 -990
rect -181 -1178 -175 -1002
rect -141 -1178 -135 -1002
rect -181 -1190 -135 -1178
rect -23 -1002 23 -990
rect -23 -1178 -17 -1002
rect 17 -1178 23 -1002
rect -23 -1190 23 -1178
rect 135 -1002 181 -990
rect 135 -1178 141 -1002
rect 175 -1178 181 -1002
rect 135 -1190 181 -1178
rect 293 -1002 339 -990
rect 293 -1178 299 -1002
rect 333 -1178 339 -1002
rect 293 -1190 339 -1178
rect 451 -1002 497 -990
rect 451 -1178 457 -1002
rect 491 -1178 497 -1002
rect 451 -1190 497 -1178
rect 609 -1002 655 -990
rect 609 -1178 615 -1002
rect 649 -1178 655 -1002
rect 609 -1190 655 -1178
rect 767 -1002 813 -990
rect 767 -1178 773 -1002
rect 807 -1178 813 -1002
rect 767 -1190 813 -1178
rect 925 -1002 971 -990
rect 925 -1178 931 -1002
rect 965 -1178 971 -1002
rect 925 -1190 971 -1178
rect 1083 -1002 1129 -990
rect 1083 -1178 1089 -1002
rect 1123 -1178 1129 -1002
rect 1083 -1190 1129 -1178
rect 1241 -1002 1287 -990
rect 1241 -1178 1247 -1002
rect 1281 -1178 1287 -1002
rect 1241 -1190 1287 -1178
rect 1399 -1002 1445 -990
rect 1399 -1178 1405 -1002
rect 1439 -1178 1445 -1002
rect 1399 -1190 1445 -1178
rect 1557 -1002 1603 -990
rect 1557 -1178 1563 -1002
rect 1597 -1178 1603 -1002
rect 1557 -1190 1603 -1178
rect -1547 -1237 -1455 -1231
rect -1547 -1271 -1535 -1237
rect -1467 -1271 -1455 -1237
rect -1547 -1277 -1455 -1271
rect -1389 -1237 -1297 -1231
rect -1389 -1271 -1377 -1237
rect -1309 -1271 -1297 -1237
rect -1389 -1277 -1297 -1271
rect -1231 -1237 -1139 -1231
rect -1231 -1271 -1219 -1237
rect -1151 -1271 -1139 -1237
rect -1231 -1277 -1139 -1271
rect -1073 -1237 -981 -1231
rect -1073 -1271 -1061 -1237
rect -993 -1271 -981 -1237
rect -1073 -1277 -981 -1271
rect -915 -1237 -823 -1231
rect -915 -1271 -903 -1237
rect -835 -1271 -823 -1237
rect -915 -1277 -823 -1271
rect -757 -1237 -665 -1231
rect -757 -1271 -745 -1237
rect -677 -1271 -665 -1237
rect -757 -1277 -665 -1271
rect -599 -1237 -507 -1231
rect -599 -1271 -587 -1237
rect -519 -1271 -507 -1237
rect -599 -1277 -507 -1271
rect -441 -1237 -349 -1231
rect -441 -1271 -429 -1237
rect -361 -1271 -349 -1237
rect -441 -1277 -349 -1271
rect -283 -1237 -191 -1231
rect -283 -1271 -271 -1237
rect -203 -1271 -191 -1237
rect -283 -1277 -191 -1271
rect -125 -1237 -33 -1231
rect -125 -1271 -113 -1237
rect -45 -1271 -33 -1237
rect -125 -1277 -33 -1271
rect 33 -1237 125 -1231
rect 33 -1271 45 -1237
rect 113 -1271 125 -1237
rect 33 -1277 125 -1271
rect 191 -1237 283 -1231
rect 191 -1271 203 -1237
rect 271 -1271 283 -1237
rect 191 -1277 283 -1271
rect 349 -1237 441 -1231
rect 349 -1271 361 -1237
rect 429 -1271 441 -1237
rect 349 -1277 441 -1271
rect 507 -1237 599 -1231
rect 507 -1271 519 -1237
rect 587 -1271 599 -1237
rect 507 -1277 599 -1271
rect 665 -1237 757 -1231
rect 665 -1271 677 -1237
rect 745 -1271 757 -1237
rect 665 -1277 757 -1271
rect 823 -1237 915 -1231
rect 823 -1271 835 -1237
rect 903 -1271 915 -1237
rect 823 -1277 915 -1271
rect 981 -1237 1073 -1231
rect 981 -1271 993 -1237
rect 1061 -1271 1073 -1237
rect 981 -1277 1073 -1271
rect 1139 -1237 1231 -1231
rect 1139 -1271 1151 -1237
rect 1219 -1271 1231 -1237
rect 1139 -1277 1231 -1271
rect 1297 -1237 1389 -1231
rect 1297 -1271 1309 -1237
rect 1377 -1271 1389 -1237
rect 1297 -1277 1389 -1271
rect 1455 -1237 1547 -1231
rect 1455 -1271 1467 -1237
rect 1535 -1271 1547 -1237
rect 1455 -1277 1547 -1271
rect -1547 -1345 -1455 -1339
rect -1547 -1379 -1535 -1345
rect -1467 -1379 -1455 -1345
rect -1547 -1385 -1455 -1379
rect -1389 -1345 -1297 -1339
rect -1389 -1379 -1377 -1345
rect -1309 -1379 -1297 -1345
rect -1389 -1385 -1297 -1379
rect -1231 -1345 -1139 -1339
rect -1231 -1379 -1219 -1345
rect -1151 -1379 -1139 -1345
rect -1231 -1385 -1139 -1379
rect -1073 -1345 -981 -1339
rect -1073 -1379 -1061 -1345
rect -993 -1379 -981 -1345
rect -1073 -1385 -981 -1379
rect -915 -1345 -823 -1339
rect -915 -1379 -903 -1345
rect -835 -1379 -823 -1345
rect -915 -1385 -823 -1379
rect -757 -1345 -665 -1339
rect -757 -1379 -745 -1345
rect -677 -1379 -665 -1345
rect -757 -1385 -665 -1379
rect -599 -1345 -507 -1339
rect -599 -1379 -587 -1345
rect -519 -1379 -507 -1345
rect -599 -1385 -507 -1379
rect -441 -1345 -349 -1339
rect -441 -1379 -429 -1345
rect -361 -1379 -349 -1345
rect -441 -1385 -349 -1379
rect -283 -1345 -191 -1339
rect -283 -1379 -271 -1345
rect -203 -1379 -191 -1345
rect -283 -1385 -191 -1379
rect -125 -1345 -33 -1339
rect -125 -1379 -113 -1345
rect -45 -1379 -33 -1345
rect -125 -1385 -33 -1379
rect 33 -1345 125 -1339
rect 33 -1379 45 -1345
rect 113 -1379 125 -1345
rect 33 -1385 125 -1379
rect 191 -1345 283 -1339
rect 191 -1379 203 -1345
rect 271 -1379 283 -1345
rect 191 -1385 283 -1379
rect 349 -1345 441 -1339
rect 349 -1379 361 -1345
rect 429 -1379 441 -1345
rect 349 -1385 441 -1379
rect 507 -1345 599 -1339
rect 507 -1379 519 -1345
rect 587 -1379 599 -1345
rect 507 -1385 599 -1379
rect 665 -1345 757 -1339
rect 665 -1379 677 -1345
rect 745 -1379 757 -1345
rect 665 -1385 757 -1379
rect 823 -1345 915 -1339
rect 823 -1379 835 -1345
rect 903 -1379 915 -1345
rect 823 -1385 915 -1379
rect 981 -1345 1073 -1339
rect 981 -1379 993 -1345
rect 1061 -1379 1073 -1345
rect 981 -1385 1073 -1379
rect 1139 -1345 1231 -1339
rect 1139 -1379 1151 -1345
rect 1219 -1379 1231 -1345
rect 1139 -1385 1231 -1379
rect 1297 -1345 1389 -1339
rect 1297 -1379 1309 -1345
rect 1377 -1379 1389 -1345
rect 1297 -1385 1389 -1379
rect 1455 -1345 1547 -1339
rect 1455 -1379 1467 -1345
rect 1535 -1379 1547 -1345
rect 1455 -1385 1547 -1379
rect -1603 -1438 -1557 -1426
rect -1603 -1614 -1597 -1438
rect -1563 -1614 -1557 -1438
rect -1603 -1626 -1557 -1614
rect -1445 -1438 -1399 -1426
rect -1445 -1614 -1439 -1438
rect -1405 -1614 -1399 -1438
rect -1445 -1626 -1399 -1614
rect -1287 -1438 -1241 -1426
rect -1287 -1614 -1281 -1438
rect -1247 -1614 -1241 -1438
rect -1287 -1626 -1241 -1614
rect -1129 -1438 -1083 -1426
rect -1129 -1614 -1123 -1438
rect -1089 -1614 -1083 -1438
rect -1129 -1626 -1083 -1614
rect -971 -1438 -925 -1426
rect -971 -1614 -965 -1438
rect -931 -1614 -925 -1438
rect -971 -1626 -925 -1614
rect -813 -1438 -767 -1426
rect -813 -1614 -807 -1438
rect -773 -1614 -767 -1438
rect -813 -1626 -767 -1614
rect -655 -1438 -609 -1426
rect -655 -1614 -649 -1438
rect -615 -1614 -609 -1438
rect -655 -1626 -609 -1614
rect -497 -1438 -451 -1426
rect -497 -1614 -491 -1438
rect -457 -1614 -451 -1438
rect -497 -1626 -451 -1614
rect -339 -1438 -293 -1426
rect -339 -1614 -333 -1438
rect -299 -1614 -293 -1438
rect -339 -1626 -293 -1614
rect -181 -1438 -135 -1426
rect -181 -1614 -175 -1438
rect -141 -1614 -135 -1438
rect -181 -1626 -135 -1614
rect -23 -1438 23 -1426
rect -23 -1614 -17 -1438
rect 17 -1614 23 -1438
rect -23 -1626 23 -1614
rect 135 -1438 181 -1426
rect 135 -1614 141 -1438
rect 175 -1614 181 -1438
rect 135 -1626 181 -1614
rect 293 -1438 339 -1426
rect 293 -1614 299 -1438
rect 333 -1614 339 -1438
rect 293 -1626 339 -1614
rect 451 -1438 497 -1426
rect 451 -1614 457 -1438
rect 491 -1614 497 -1438
rect 451 -1626 497 -1614
rect 609 -1438 655 -1426
rect 609 -1614 615 -1438
rect 649 -1614 655 -1438
rect 609 -1626 655 -1614
rect 767 -1438 813 -1426
rect 767 -1614 773 -1438
rect 807 -1614 813 -1438
rect 767 -1626 813 -1614
rect 925 -1438 971 -1426
rect 925 -1614 931 -1438
rect 965 -1614 971 -1438
rect 925 -1626 971 -1614
rect 1083 -1438 1129 -1426
rect 1083 -1614 1089 -1438
rect 1123 -1614 1129 -1438
rect 1083 -1626 1129 -1614
rect 1241 -1438 1287 -1426
rect 1241 -1614 1247 -1438
rect 1281 -1614 1287 -1438
rect 1241 -1626 1287 -1614
rect 1399 -1438 1445 -1426
rect 1399 -1614 1405 -1438
rect 1439 -1614 1445 -1438
rect 1399 -1626 1445 -1614
rect 1557 -1438 1603 -1426
rect 1557 -1614 1563 -1438
rect 1597 -1614 1603 -1438
rect 1557 -1626 1603 -1614
rect -1547 -1673 -1455 -1667
rect -1547 -1707 -1535 -1673
rect -1467 -1707 -1455 -1673
rect -1547 -1713 -1455 -1707
rect -1389 -1673 -1297 -1667
rect -1389 -1707 -1377 -1673
rect -1309 -1707 -1297 -1673
rect -1389 -1713 -1297 -1707
rect -1231 -1673 -1139 -1667
rect -1231 -1707 -1219 -1673
rect -1151 -1707 -1139 -1673
rect -1231 -1713 -1139 -1707
rect -1073 -1673 -981 -1667
rect -1073 -1707 -1061 -1673
rect -993 -1707 -981 -1673
rect -1073 -1713 -981 -1707
rect -915 -1673 -823 -1667
rect -915 -1707 -903 -1673
rect -835 -1707 -823 -1673
rect -915 -1713 -823 -1707
rect -757 -1673 -665 -1667
rect -757 -1707 -745 -1673
rect -677 -1707 -665 -1673
rect -757 -1713 -665 -1707
rect -599 -1673 -507 -1667
rect -599 -1707 -587 -1673
rect -519 -1707 -507 -1673
rect -599 -1713 -507 -1707
rect -441 -1673 -349 -1667
rect -441 -1707 -429 -1673
rect -361 -1707 -349 -1673
rect -441 -1713 -349 -1707
rect -283 -1673 -191 -1667
rect -283 -1707 -271 -1673
rect -203 -1707 -191 -1673
rect -283 -1713 -191 -1707
rect -125 -1673 -33 -1667
rect -125 -1707 -113 -1673
rect -45 -1707 -33 -1673
rect -125 -1713 -33 -1707
rect 33 -1673 125 -1667
rect 33 -1707 45 -1673
rect 113 -1707 125 -1673
rect 33 -1713 125 -1707
rect 191 -1673 283 -1667
rect 191 -1707 203 -1673
rect 271 -1707 283 -1673
rect 191 -1713 283 -1707
rect 349 -1673 441 -1667
rect 349 -1707 361 -1673
rect 429 -1707 441 -1673
rect 349 -1713 441 -1707
rect 507 -1673 599 -1667
rect 507 -1707 519 -1673
rect 587 -1707 599 -1673
rect 507 -1713 599 -1707
rect 665 -1673 757 -1667
rect 665 -1707 677 -1673
rect 745 -1707 757 -1673
rect 665 -1713 757 -1707
rect 823 -1673 915 -1667
rect 823 -1707 835 -1673
rect 903 -1707 915 -1673
rect 823 -1713 915 -1707
rect 981 -1673 1073 -1667
rect 981 -1707 993 -1673
rect 1061 -1707 1073 -1673
rect 981 -1713 1073 -1707
rect 1139 -1673 1231 -1667
rect 1139 -1707 1151 -1673
rect 1219 -1707 1231 -1673
rect 1139 -1713 1231 -1707
rect 1297 -1673 1389 -1667
rect 1297 -1707 1309 -1673
rect 1377 -1707 1389 -1673
rect 1297 -1713 1389 -1707
rect 1455 -1673 1547 -1667
rect 1455 -1707 1467 -1673
rect 1535 -1707 1547 -1673
rect 1455 -1713 1547 -1707
rect -1547 -1781 -1455 -1775
rect -1547 -1815 -1535 -1781
rect -1467 -1815 -1455 -1781
rect -1547 -1821 -1455 -1815
rect -1389 -1781 -1297 -1775
rect -1389 -1815 -1377 -1781
rect -1309 -1815 -1297 -1781
rect -1389 -1821 -1297 -1815
rect -1231 -1781 -1139 -1775
rect -1231 -1815 -1219 -1781
rect -1151 -1815 -1139 -1781
rect -1231 -1821 -1139 -1815
rect -1073 -1781 -981 -1775
rect -1073 -1815 -1061 -1781
rect -993 -1815 -981 -1781
rect -1073 -1821 -981 -1815
rect -915 -1781 -823 -1775
rect -915 -1815 -903 -1781
rect -835 -1815 -823 -1781
rect -915 -1821 -823 -1815
rect -757 -1781 -665 -1775
rect -757 -1815 -745 -1781
rect -677 -1815 -665 -1781
rect -757 -1821 -665 -1815
rect -599 -1781 -507 -1775
rect -599 -1815 -587 -1781
rect -519 -1815 -507 -1781
rect -599 -1821 -507 -1815
rect -441 -1781 -349 -1775
rect -441 -1815 -429 -1781
rect -361 -1815 -349 -1781
rect -441 -1821 -349 -1815
rect -283 -1781 -191 -1775
rect -283 -1815 -271 -1781
rect -203 -1815 -191 -1781
rect -283 -1821 -191 -1815
rect -125 -1781 -33 -1775
rect -125 -1815 -113 -1781
rect -45 -1815 -33 -1781
rect -125 -1821 -33 -1815
rect 33 -1781 125 -1775
rect 33 -1815 45 -1781
rect 113 -1815 125 -1781
rect 33 -1821 125 -1815
rect 191 -1781 283 -1775
rect 191 -1815 203 -1781
rect 271 -1815 283 -1781
rect 191 -1821 283 -1815
rect 349 -1781 441 -1775
rect 349 -1815 361 -1781
rect 429 -1815 441 -1781
rect 349 -1821 441 -1815
rect 507 -1781 599 -1775
rect 507 -1815 519 -1781
rect 587 -1815 599 -1781
rect 507 -1821 599 -1815
rect 665 -1781 757 -1775
rect 665 -1815 677 -1781
rect 745 -1815 757 -1781
rect 665 -1821 757 -1815
rect 823 -1781 915 -1775
rect 823 -1815 835 -1781
rect 903 -1815 915 -1781
rect 823 -1821 915 -1815
rect 981 -1781 1073 -1775
rect 981 -1815 993 -1781
rect 1061 -1815 1073 -1781
rect 981 -1821 1073 -1815
rect 1139 -1781 1231 -1775
rect 1139 -1815 1151 -1781
rect 1219 -1815 1231 -1781
rect 1139 -1821 1231 -1815
rect 1297 -1781 1389 -1775
rect 1297 -1815 1309 -1781
rect 1377 -1815 1389 -1781
rect 1297 -1821 1389 -1815
rect 1455 -1781 1547 -1775
rect 1455 -1815 1467 -1781
rect 1535 -1815 1547 -1781
rect 1455 -1821 1547 -1815
rect -1603 -1874 -1557 -1862
rect -1603 -2050 -1597 -1874
rect -1563 -2050 -1557 -1874
rect -1603 -2062 -1557 -2050
rect -1445 -1874 -1399 -1862
rect -1445 -2050 -1439 -1874
rect -1405 -2050 -1399 -1874
rect -1445 -2062 -1399 -2050
rect -1287 -1874 -1241 -1862
rect -1287 -2050 -1281 -1874
rect -1247 -2050 -1241 -1874
rect -1287 -2062 -1241 -2050
rect -1129 -1874 -1083 -1862
rect -1129 -2050 -1123 -1874
rect -1089 -2050 -1083 -1874
rect -1129 -2062 -1083 -2050
rect -971 -1874 -925 -1862
rect -971 -2050 -965 -1874
rect -931 -2050 -925 -1874
rect -971 -2062 -925 -2050
rect -813 -1874 -767 -1862
rect -813 -2050 -807 -1874
rect -773 -2050 -767 -1874
rect -813 -2062 -767 -2050
rect -655 -1874 -609 -1862
rect -655 -2050 -649 -1874
rect -615 -2050 -609 -1874
rect -655 -2062 -609 -2050
rect -497 -1874 -451 -1862
rect -497 -2050 -491 -1874
rect -457 -2050 -451 -1874
rect -497 -2062 -451 -2050
rect -339 -1874 -293 -1862
rect -339 -2050 -333 -1874
rect -299 -2050 -293 -1874
rect -339 -2062 -293 -2050
rect -181 -1874 -135 -1862
rect -181 -2050 -175 -1874
rect -141 -2050 -135 -1874
rect -181 -2062 -135 -2050
rect -23 -1874 23 -1862
rect -23 -2050 -17 -1874
rect 17 -2050 23 -1874
rect -23 -2062 23 -2050
rect 135 -1874 181 -1862
rect 135 -2050 141 -1874
rect 175 -2050 181 -1874
rect 135 -2062 181 -2050
rect 293 -1874 339 -1862
rect 293 -2050 299 -1874
rect 333 -2050 339 -1874
rect 293 -2062 339 -2050
rect 451 -1874 497 -1862
rect 451 -2050 457 -1874
rect 491 -2050 497 -1874
rect 451 -2062 497 -2050
rect 609 -1874 655 -1862
rect 609 -2050 615 -1874
rect 649 -2050 655 -1874
rect 609 -2062 655 -2050
rect 767 -1874 813 -1862
rect 767 -2050 773 -1874
rect 807 -2050 813 -1874
rect 767 -2062 813 -2050
rect 925 -1874 971 -1862
rect 925 -2050 931 -1874
rect 965 -2050 971 -1874
rect 925 -2062 971 -2050
rect 1083 -1874 1129 -1862
rect 1083 -2050 1089 -1874
rect 1123 -2050 1129 -1874
rect 1083 -2062 1129 -2050
rect 1241 -1874 1287 -1862
rect 1241 -2050 1247 -1874
rect 1281 -2050 1287 -1874
rect 1241 -2062 1287 -2050
rect 1399 -1874 1445 -1862
rect 1399 -2050 1405 -1874
rect 1439 -2050 1445 -1874
rect 1399 -2062 1445 -2050
rect 1557 -1874 1603 -1862
rect 1557 -2050 1563 -1874
rect 1597 -2050 1603 -1874
rect 1557 -2062 1603 -2050
rect -1547 -2109 -1455 -2103
rect -1547 -2143 -1535 -2109
rect -1467 -2143 -1455 -2109
rect -1547 -2149 -1455 -2143
rect -1389 -2109 -1297 -2103
rect -1389 -2143 -1377 -2109
rect -1309 -2143 -1297 -2109
rect -1389 -2149 -1297 -2143
rect -1231 -2109 -1139 -2103
rect -1231 -2143 -1219 -2109
rect -1151 -2143 -1139 -2109
rect -1231 -2149 -1139 -2143
rect -1073 -2109 -981 -2103
rect -1073 -2143 -1061 -2109
rect -993 -2143 -981 -2109
rect -1073 -2149 -981 -2143
rect -915 -2109 -823 -2103
rect -915 -2143 -903 -2109
rect -835 -2143 -823 -2109
rect -915 -2149 -823 -2143
rect -757 -2109 -665 -2103
rect -757 -2143 -745 -2109
rect -677 -2143 -665 -2109
rect -757 -2149 -665 -2143
rect -599 -2109 -507 -2103
rect -599 -2143 -587 -2109
rect -519 -2143 -507 -2109
rect -599 -2149 -507 -2143
rect -441 -2109 -349 -2103
rect -441 -2143 -429 -2109
rect -361 -2143 -349 -2109
rect -441 -2149 -349 -2143
rect -283 -2109 -191 -2103
rect -283 -2143 -271 -2109
rect -203 -2143 -191 -2109
rect -283 -2149 -191 -2143
rect -125 -2109 -33 -2103
rect -125 -2143 -113 -2109
rect -45 -2143 -33 -2109
rect -125 -2149 -33 -2143
rect 33 -2109 125 -2103
rect 33 -2143 45 -2109
rect 113 -2143 125 -2109
rect 33 -2149 125 -2143
rect 191 -2109 283 -2103
rect 191 -2143 203 -2109
rect 271 -2143 283 -2109
rect 191 -2149 283 -2143
rect 349 -2109 441 -2103
rect 349 -2143 361 -2109
rect 429 -2143 441 -2109
rect 349 -2149 441 -2143
rect 507 -2109 599 -2103
rect 507 -2143 519 -2109
rect 587 -2143 599 -2109
rect 507 -2149 599 -2143
rect 665 -2109 757 -2103
rect 665 -2143 677 -2109
rect 745 -2143 757 -2109
rect 665 -2149 757 -2143
rect 823 -2109 915 -2103
rect 823 -2143 835 -2109
rect 903 -2143 915 -2109
rect 823 -2149 915 -2143
rect 981 -2109 1073 -2103
rect 981 -2143 993 -2109
rect 1061 -2143 1073 -2109
rect 981 -2149 1073 -2143
rect 1139 -2109 1231 -2103
rect 1139 -2143 1151 -2109
rect 1219 -2143 1231 -2109
rect 1139 -2149 1231 -2143
rect 1297 -2109 1389 -2103
rect 1297 -2143 1309 -2109
rect 1377 -2143 1389 -2109
rect 1297 -2149 1389 -2143
rect 1455 -2109 1547 -2103
rect 1455 -2143 1467 -2109
rect 1535 -2143 1547 -2109
rect 1455 -2149 1547 -2143
rect -1547 -2217 -1455 -2211
rect -1547 -2251 -1535 -2217
rect -1467 -2251 -1455 -2217
rect -1547 -2257 -1455 -2251
rect -1389 -2217 -1297 -2211
rect -1389 -2251 -1377 -2217
rect -1309 -2251 -1297 -2217
rect -1389 -2257 -1297 -2251
rect -1231 -2217 -1139 -2211
rect -1231 -2251 -1219 -2217
rect -1151 -2251 -1139 -2217
rect -1231 -2257 -1139 -2251
rect -1073 -2217 -981 -2211
rect -1073 -2251 -1061 -2217
rect -993 -2251 -981 -2217
rect -1073 -2257 -981 -2251
rect -915 -2217 -823 -2211
rect -915 -2251 -903 -2217
rect -835 -2251 -823 -2217
rect -915 -2257 -823 -2251
rect -757 -2217 -665 -2211
rect -757 -2251 -745 -2217
rect -677 -2251 -665 -2217
rect -757 -2257 -665 -2251
rect -599 -2217 -507 -2211
rect -599 -2251 -587 -2217
rect -519 -2251 -507 -2217
rect -599 -2257 -507 -2251
rect -441 -2217 -349 -2211
rect -441 -2251 -429 -2217
rect -361 -2251 -349 -2217
rect -441 -2257 -349 -2251
rect -283 -2217 -191 -2211
rect -283 -2251 -271 -2217
rect -203 -2251 -191 -2217
rect -283 -2257 -191 -2251
rect -125 -2217 -33 -2211
rect -125 -2251 -113 -2217
rect -45 -2251 -33 -2217
rect -125 -2257 -33 -2251
rect 33 -2217 125 -2211
rect 33 -2251 45 -2217
rect 113 -2251 125 -2217
rect 33 -2257 125 -2251
rect 191 -2217 283 -2211
rect 191 -2251 203 -2217
rect 271 -2251 283 -2217
rect 191 -2257 283 -2251
rect 349 -2217 441 -2211
rect 349 -2251 361 -2217
rect 429 -2251 441 -2217
rect 349 -2257 441 -2251
rect 507 -2217 599 -2211
rect 507 -2251 519 -2217
rect 587 -2251 599 -2217
rect 507 -2257 599 -2251
rect 665 -2217 757 -2211
rect 665 -2251 677 -2217
rect 745 -2251 757 -2217
rect 665 -2257 757 -2251
rect 823 -2217 915 -2211
rect 823 -2251 835 -2217
rect 903 -2251 915 -2217
rect 823 -2257 915 -2251
rect 981 -2217 1073 -2211
rect 981 -2251 993 -2217
rect 1061 -2251 1073 -2217
rect 981 -2257 1073 -2251
rect 1139 -2217 1231 -2211
rect 1139 -2251 1151 -2217
rect 1219 -2251 1231 -2217
rect 1139 -2257 1231 -2251
rect 1297 -2217 1389 -2211
rect 1297 -2251 1309 -2217
rect 1377 -2251 1389 -2217
rect 1297 -2257 1389 -2251
rect 1455 -2217 1547 -2211
rect 1455 -2251 1467 -2217
rect 1535 -2251 1547 -2217
rect 1455 -2257 1547 -2251
rect -1603 -2310 -1557 -2298
rect -1603 -2486 -1597 -2310
rect -1563 -2486 -1557 -2310
rect -1603 -2498 -1557 -2486
rect -1445 -2310 -1399 -2298
rect -1445 -2486 -1439 -2310
rect -1405 -2486 -1399 -2310
rect -1445 -2498 -1399 -2486
rect -1287 -2310 -1241 -2298
rect -1287 -2486 -1281 -2310
rect -1247 -2486 -1241 -2310
rect -1287 -2498 -1241 -2486
rect -1129 -2310 -1083 -2298
rect -1129 -2486 -1123 -2310
rect -1089 -2486 -1083 -2310
rect -1129 -2498 -1083 -2486
rect -971 -2310 -925 -2298
rect -971 -2486 -965 -2310
rect -931 -2486 -925 -2310
rect -971 -2498 -925 -2486
rect -813 -2310 -767 -2298
rect -813 -2486 -807 -2310
rect -773 -2486 -767 -2310
rect -813 -2498 -767 -2486
rect -655 -2310 -609 -2298
rect -655 -2486 -649 -2310
rect -615 -2486 -609 -2310
rect -655 -2498 -609 -2486
rect -497 -2310 -451 -2298
rect -497 -2486 -491 -2310
rect -457 -2486 -451 -2310
rect -497 -2498 -451 -2486
rect -339 -2310 -293 -2298
rect -339 -2486 -333 -2310
rect -299 -2486 -293 -2310
rect -339 -2498 -293 -2486
rect -181 -2310 -135 -2298
rect -181 -2486 -175 -2310
rect -141 -2486 -135 -2310
rect -181 -2498 -135 -2486
rect -23 -2310 23 -2298
rect -23 -2486 -17 -2310
rect 17 -2486 23 -2310
rect -23 -2498 23 -2486
rect 135 -2310 181 -2298
rect 135 -2486 141 -2310
rect 175 -2486 181 -2310
rect 135 -2498 181 -2486
rect 293 -2310 339 -2298
rect 293 -2486 299 -2310
rect 333 -2486 339 -2310
rect 293 -2498 339 -2486
rect 451 -2310 497 -2298
rect 451 -2486 457 -2310
rect 491 -2486 497 -2310
rect 451 -2498 497 -2486
rect 609 -2310 655 -2298
rect 609 -2486 615 -2310
rect 649 -2486 655 -2310
rect 609 -2498 655 -2486
rect 767 -2310 813 -2298
rect 767 -2486 773 -2310
rect 807 -2486 813 -2310
rect 767 -2498 813 -2486
rect 925 -2310 971 -2298
rect 925 -2486 931 -2310
rect 965 -2486 971 -2310
rect 925 -2498 971 -2486
rect 1083 -2310 1129 -2298
rect 1083 -2486 1089 -2310
rect 1123 -2486 1129 -2310
rect 1083 -2498 1129 -2486
rect 1241 -2310 1287 -2298
rect 1241 -2486 1247 -2310
rect 1281 -2486 1287 -2310
rect 1241 -2498 1287 -2486
rect 1399 -2310 1445 -2298
rect 1399 -2486 1405 -2310
rect 1439 -2486 1445 -2310
rect 1399 -2498 1445 -2486
rect 1557 -2310 1603 -2298
rect 1557 -2486 1563 -2310
rect 1597 -2486 1603 -2310
rect 1557 -2498 1603 -2486
rect -1547 -2545 -1455 -2539
rect -1547 -2579 -1535 -2545
rect -1467 -2579 -1455 -2545
rect -1547 -2585 -1455 -2579
rect -1389 -2545 -1297 -2539
rect -1389 -2579 -1377 -2545
rect -1309 -2579 -1297 -2545
rect -1389 -2585 -1297 -2579
rect -1231 -2545 -1139 -2539
rect -1231 -2579 -1219 -2545
rect -1151 -2579 -1139 -2545
rect -1231 -2585 -1139 -2579
rect -1073 -2545 -981 -2539
rect -1073 -2579 -1061 -2545
rect -993 -2579 -981 -2545
rect -1073 -2585 -981 -2579
rect -915 -2545 -823 -2539
rect -915 -2579 -903 -2545
rect -835 -2579 -823 -2545
rect -915 -2585 -823 -2579
rect -757 -2545 -665 -2539
rect -757 -2579 -745 -2545
rect -677 -2579 -665 -2545
rect -757 -2585 -665 -2579
rect -599 -2545 -507 -2539
rect -599 -2579 -587 -2545
rect -519 -2579 -507 -2545
rect -599 -2585 -507 -2579
rect -441 -2545 -349 -2539
rect -441 -2579 -429 -2545
rect -361 -2579 -349 -2545
rect -441 -2585 -349 -2579
rect -283 -2545 -191 -2539
rect -283 -2579 -271 -2545
rect -203 -2579 -191 -2545
rect -283 -2585 -191 -2579
rect -125 -2545 -33 -2539
rect -125 -2579 -113 -2545
rect -45 -2579 -33 -2545
rect -125 -2585 -33 -2579
rect 33 -2545 125 -2539
rect 33 -2579 45 -2545
rect 113 -2579 125 -2545
rect 33 -2585 125 -2579
rect 191 -2545 283 -2539
rect 191 -2579 203 -2545
rect 271 -2579 283 -2545
rect 191 -2585 283 -2579
rect 349 -2545 441 -2539
rect 349 -2579 361 -2545
rect 429 -2579 441 -2545
rect 349 -2585 441 -2579
rect 507 -2545 599 -2539
rect 507 -2579 519 -2545
rect 587 -2579 599 -2545
rect 507 -2585 599 -2579
rect 665 -2545 757 -2539
rect 665 -2579 677 -2545
rect 745 -2579 757 -2545
rect 665 -2585 757 -2579
rect 823 -2545 915 -2539
rect 823 -2579 835 -2545
rect 903 -2579 915 -2545
rect 823 -2585 915 -2579
rect 981 -2545 1073 -2539
rect 981 -2579 993 -2545
rect 1061 -2579 1073 -2545
rect 981 -2585 1073 -2579
rect 1139 -2545 1231 -2539
rect 1139 -2579 1151 -2545
rect 1219 -2579 1231 -2545
rect 1139 -2585 1231 -2579
rect 1297 -2545 1389 -2539
rect 1297 -2579 1309 -2545
rect 1377 -2579 1389 -2545
rect 1297 -2585 1389 -2579
rect 1455 -2545 1547 -2539
rect 1455 -2579 1467 -2545
rect 1535 -2579 1547 -2545
rect 1455 -2585 1547 -2579
rect -1547 -2653 -1455 -2647
rect -1547 -2687 -1535 -2653
rect -1467 -2687 -1455 -2653
rect -1547 -2693 -1455 -2687
rect -1389 -2653 -1297 -2647
rect -1389 -2687 -1377 -2653
rect -1309 -2687 -1297 -2653
rect -1389 -2693 -1297 -2687
rect -1231 -2653 -1139 -2647
rect -1231 -2687 -1219 -2653
rect -1151 -2687 -1139 -2653
rect -1231 -2693 -1139 -2687
rect -1073 -2653 -981 -2647
rect -1073 -2687 -1061 -2653
rect -993 -2687 -981 -2653
rect -1073 -2693 -981 -2687
rect -915 -2653 -823 -2647
rect -915 -2687 -903 -2653
rect -835 -2687 -823 -2653
rect -915 -2693 -823 -2687
rect -757 -2653 -665 -2647
rect -757 -2687 -745 -2653
rect -677 -2687 -665 -2653
rect -757 -2693 -665 -2687
rect -599 -2653 -507 -2647
rect -599 -2687 -587 -2653
rect -519 -2687 -507 -2653
rect -599 -2693 -507 -2687
rect -441 -2653 -349 -2647
rect -441 -2687 -429 -2653
rect -361 -2687 -349 -2653
rect -441 -2693 -349 -2687
rect -283 -2653 -191 -2647
rect -283 -2687 -271 -2653
rect -203 -2687 -191 -2653
rect -283 -2693 -191 -2687
rect -125 -2653 -33 -2647
rect -125 -2687 -113 -2653
rect -45 -2687 -33 -2653
rect -125 -2693 -33 -2687
rect 33 -2653 125 -2647
rect 33 -2687 45 -2653
rect 113 -2687 125 -2653
rect 33 -2693 125 -2687
rect 191 -2653 283 -2647
rect 191 -2687 203 -2653
rect 271 -2687 283 -2653
rect 191 -2693 283 -2687
rect 349 -2653 441 -2647
rect 349 -2687 361 -2653
rect 429 -2687 441 -2653
rect 349 -2693 441 -2687
rect 507 -2653 599 -2647
rect 507 -2687 519 -2653
rect 587 -2687 599 -2653
rect 507 -2693 599 -2687
rect 665 -2653 757 -2647
rect 665 -2687 677 -2653
rect 745 -2687 757 -2653
rect 665 -2693 757 -2687
rect 823 -2653 915 -2647
rect 823 -2687 835 -2653
rect 903 -2687 915 -2653
rect 823 -2693 915 -2687
rect 981 -2653 1073 -2647
rect 981 -2687 993 -2653
rect 1061 -2687 1073 -2653
rect 981 -2693 1073 -2687
rect 1139 -2653 1231 -2647
rect 1139 -2687 1151 -2653
rect 1219 -2687 1231 -2653
rect 1139 -2693 1231 -2687
rect 1297 -2653 1389 -2647
rect 1297 -2687 1309 -2653
rect 1377 -2687 1389 -2653
rect 1297 -2693 1389 -2687
rect 1455 -2653 1547 -2647
rect 1455 -2687 1467 -2653
rect 1535 -2687 1547 -2653
rect 1455 -2693 1547 -2687
rect -1603 -2746 -1557 -2734
rect -1603 -2922 -1597 -2746
rect -1563 -2922 -1557 -2746
rect -1603 -2934 -1557 -2922
rect -1445 -2746 -1399 -2734
rect -1445 -2922 -1439 -2746
rect -1405 -2922 -1399 -2746
rect -1445 -2934 -1399 -2922
rect -1287 -2746 -1241 -2734
rect -1287 -2922 -1281 -2746
rect -1247 -2922 -1241 -2746
rect -1287 -2934 -1241 -2922
rect -1129 -2746 -1083 -2734
rect -1129 -2922 -1123 -2746
rect -1089 -2922 -1083 -2746
rect -1129 -2934 -1083 -2922
rect -971 -2746 -925 -2734
rect -971 -2922 -965 -2746
rect -931 -2922 -925 -2746
rect -971 -2934 -925 -2922
rect -813 -2746 -767 -2734
rect -813 -2922 -807 -2746
rect -773 -2922 -767 -2746
rect -813 -2934 -767 -2922
rect -655 -2746 -609 -2734
rect -655 -2922 -649 -2746
rect -615 -2922 -609 -2746
rect -655 -2934 -609 -2922
rect -497 -2746 -451 -2734
rect -497 -2922 -491 -2746
rect -457 -2922 -451 -2746
rect -497 -2934 -451 -2922
rect -339 -2746 -293 -2734
rect -339 -2922 -333 -2746
rect -299 -2922 -293 -2746
rect -339 -2934 -293 -2922
rect -181 -2746 -135 -2734
rect -181 -2922 -175 -2746
rect -141 -2922 -135 -2746
rect -181 -2934 -135 -2922
rect -23 -2746 23 -2734
rect -23 -2922 -17 -2746
rect 17 -2922 23 -2746
rect -23 -2934 23 -2922
rect 135 -2746 181 -2734
rect 135 -2922 141 -2746
rect 175 -2922 181 -2746
rect 135 -2934 181 -2922
rect 293 -2746 339 -2734
rect 293 -2922 299 -2746
rect 333 -2922 339 -2746
rect 293 -2934 339 -2922
rect 451 -2746 497 -2734
rect 451 -2922 457 -2746
rect 491 -2922 497 -2746
rect 451 -2934 497 -2922
rect 609 -2746 655 -2734
rect 609 -2922 615 -2746
rect 649 -2922 655 -2746
rect 609 -2934 655 -2922
rect 767 -2746 813 -2734
rect 767 -2922 773 -2746
rect 807 -2922 813 -2746
rect 767 -2934 813 -2922
rect 925 -2746 971 -2734
rect 925 -2922 931 -2746
rect 965 -2922 971 -2746
rect 925 -2934 971 -2922
rect 1083 -2746 1129 -2734
rect 1083 -2922 1089 -2746
rect 1123 -2922 1129 -2746
rect 1083 -2934 1129 -2922
rect 1241 -2746 1287 -2734
rect 1241 -2922 1247 -2746
rect 1281 -2922 1287 -2746
rect 1241 -2934 1287 -2922
rect 1399 -2746 1445 -2734
rect 1399 -2922 1405 -2746
rect 1439 -2922 1445 -2746
rect 1399 -2934 1445 -2922
rect 1557 -2746 1603 -2734
rect 1557 -2922 1563 -2746
rect 1597 -2922 1603 -2746
rect 1557 -2934 1603 -2922
rect -1547 -2981 -1455 -2975
rect -1547 -3015 -1535 -2981
rect -1467 -3015 -1455 -2981
rect -1547 -3021 -1455 -3015
rect -1389 -2981 -1297 -2975
rect -1389 -3015 -1377 -2981
rect -1309 -3015 -1297 -2981
rect -1389 -3021 -1297 -3015
rect -1231 -2981 -1139 -2975
rect -1231 -3015 -1219 -2981
rect -1151 -3015 -1139 -2981
rect -1231 -3021 -1139 -3015
rect -1073 -2981 -981 -2975
rect -1073 -3015 -1061 -2981
rect -993 -3015 -981 -2981
rect -1073 -3021 -981 -3015
rect -915 -2981 -823 -2975
rect -915 -3015 -903 -2981
rect -835 -3015 -823 -2981
rect -915 -3021 -823 -3015
rect -757 -2981 -665 -2975
rect -757 -3015 -745 -2981
rect -677 -3015 -665 -2981
rect -757 -3021 -665 -3015
rect -599 -2981 -507 -2975
rect -599 -3015 -587 -2981
rect -519 -3015 -507 -2981
rect -599 -3021 -507 -3015
rect -441 -2981 -349 -2975
rect -441 -3015 -429 -2981
rect -361 -3015 -349 -2981
rect -441 -3021 -349 -3015
rect -283 -2981 -191 -2975
rect -283 -3015 -271 -2981
rect -203 -3015 -191 -2981
rect -283 -3021 -191 -3015
rect -125 -2981 -33 -2975
rect -125 -3015 -113 -2981
rect -45 -3015 -33 -2981
rect -125 -3021 -33 -3015
rect 33 -2981 125 -2975
rect 33 -3015 45 -2981
rect 113 -3015 125 -2981
rect 33 -3021 125 -3015
rect 191 -2981 283 -2975
rect 191 -3015 203 -2981
rect 271 -3015 283 -2981
rect 191 -3021 283 -3015
rect 349 -2981 441 -2975
rect 349 -3015 361 -2981
rect 429 -3015 441 -2981
rect 349 -3021 441 -3015
rect 507 -2981 599 -2975
rect 507 -3015 519 -2981
rect 587 -3015 599 -2981
rect 507 -3021 599 -3015
rect 665 -2981 757 -2975
rect 665 -3015 677 -2981
rect 745 -3015 757 -2981
rect 665 -3021 757 -3015
rect 823 -2981 915 -2975
rect 823 -3015 835 -2981
rect 903 -3015 915 -2981
rect 823 -3021 915 -3015
rect 981 -2981 1073 -2975
rect 981 -3015 993 -2981
rect 1061 -3015 1073 -2981
rect 981 -3021 1073 -3015
rect 1139 -2981 1231 -2975
rect 1139 -3015 1151 -2981
rect 1219 -3015 1231 -2981
rect 1139 -3021 1231 -3015
rect 1297 -2981 1389 -2975
rect 1297 -3015 1309 -2981
rect 1377 -3015 1389 -2981
rect 1297 -3021 1389 -3015
rect 1455 -2981 1547 -2975
rect 1455 -3015 1467 -2981
rect 1535 -3015 1547 -2981
rect 1455 -3021 1547 -3015
<< properties >>
string FIXED_BBOX -1714 -3136 1714 3136
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.5 m 14 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
