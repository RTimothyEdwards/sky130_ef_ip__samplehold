magic
tech sky130A
magscale 1 2
timestamp 1718244471
<< locali >>
rect 1350 10646 1667 10669
rect 1350 10489 1373 10646
rect 1642 10489 1667 10646
rect 1350 10454 1667 10489
rect 1475 9831 1605 10454
rect 1094 9512 1374 9534
rect 1094 9423 1112 9512
rect 1355 9423 1374 9512
rect 1094 9400 1374 9423
rect 2935 8813 3044 8842
rect 2935 8404 2951 8813
rect 3020 8404 3044 8813
rect 2935 8380 3044 8404
rect 2938 7988 3041 8016
rect 2938 7579 2955 7988
rect 3024 7579 3041 7988
rect 2938 7555 3041 7579
rect 1094 7000 1374 7024
rect 1094 6911 1113 7000
rect 1356 6911 1374 7000
rect 1094 6890 1374 6911
rect 1512 6154 1642 6597
rect 1351 6116 1668 6154
rect 1351 5904 1378 6116
rect 1635 5904 1668 6116
rect 1351 5877 1668 5904
<< viali >>
rect 1373 10489 1642 10646
rect 1112 9423 1355 9512
rect 2951 8404 3020 8813
rect 2955 7579 3024 7988
rect 1113 6911 1356 7000
rect 1378 5904 1635 6116
<< metal1 >>
rect 671 11512 14883 11558
rect 671 11264 14397 11512
rect 671 10817 2263 11264
rect 2775 10841 14397 11264
rect 14842 10841 14883 11512
rect 2775 10817 14883 10841
rect 671 10797 14883 10817
rect 1350 10646 3811 10670
rect 1350 10489 1373 10646
rect 1642 10563 3811 10646
rect 1642 10489 1667 10563
rect 1350 10454 1667 10489
rect 3300 10327 3642 10349
rect 1322 10016 1368 10317
rect 778 9970 1368 10016
rect 3300 10009 3320 10327
rect 3623 10009 3642 10327
rect 778 9558 824 9970
rect 875 9848 2996 9850
rect 875 9741 1368 9848
rect 1659 9741 2996 9848
rect 589 9500 824 9558
rect 1094 9512 1374 9534
rect 1094 9500 1112 9512
rect 589 9431 1112 9500
rect 589 9358 786 9431
rect 1094 9423 1112 9431
rect 1355 9423 1374 9512
rect 1094 9400 1374 9423
rect 3300 9151 3642 10009
rect 678 9137 1225 9151
rect 2970 9137 3642 9151
rect 678 9127 3642 9137
rect 678 8867 704 9127
rect 1200 8921 3642 9127
rect 1200 8867 1225 8921
rect 2970 8901 3642 8921
rect 678 8842 1225 8867
rect 2935 8813 3044 8842
rect 2935 8404 2951 8813
rect 3020 8430 3044 8813
rect 3020 8404 3188 8430
rect 2935 8380 3188 8404
rect 2982 8379 3188 8380
rect 874 8304 2982 8313
rect 874 8099 1368 8304
rect 1650 8099 2982 8304
rect 874 8097 2982 8099
rect 2938 7988 3087 8016
rect 685 7565 1226 7595
rect 685 7300 708 7565
rect 1199 7511 1226 7565
rect 2938 7579 2955 7988
rect 3024 7579 3087 7988
rect 2938 7555 3087 7579
rect 1199 7300 2985 7511
rect 685 7295 2985 7300
rect 685 7276 1226 7295
rect 1800 7244 2118 7245
rect 1800 7170 1808 7244
rect 2108 7170 2118 7244
rect 1800 7158 2118 7170
rect 589 6989 789 7042
rect 1094 7000 1374 7024
rect 1094 6989 1113 7000
rect 589 6920 1113 6989
rect 589 6842 824 6920
rect 1094 6911 1113 6920
rect 1356 6911 1374 7000
rect 1094 6890 1374 6911
rect 775 6443 824 6842
rect 878 6565 1364 6696
rect 1660 6565 2984 6696
rect 878 6563 2984 6565
rect 2264 6454 2759 6496
rect 775 6394 1392 6443
rect 1343 6229 1392 6394
rect 1351 6154 1392 6155
rect 1351 6116 1668 6154
rect 1351 5904 1378 6116
rect 1635 5904 1668 6116
rect 2264 6126 2309 6454
rect 2715 6126 2759 6454
rect 2264 5948 2759 6126
rect 1351 5877 1668 5904
rect 2262 5937 2759 5948
rect 2262 5670 2758 5937
rect 3038 5476 3087 7555
rect 3137 6859 3188 8379
rect 3137 6760 3191 6859
rect 3137 5456 3188 6760
rect 3300 6169 3642 8901
rect 3300 6136 14803 6169
rect 3300 5555 7191 6136
rect 7795 5589 10413 6136
rect 11027 6122 14803 6136
rect 11027 5589 13849 6122
rect 7795 5575 13849 5589
rect 14463 5575 14803 6122
rect 7795 5555 14803 5575
rect 3300 5527 14803 5555
rect 2730 3979 3443 4179
rect 3643 3979 3650 4179
rect 704 2862 1160 2891
rect 704 2141 738 2862
rect 1127 2141 1160 2862
rect 704 2099 1160 2141
rect 2709 1924 3041 1994
rect 2865 1198 3218 1217
rect 2865 1012 2877 1198
rect 3204 1155 3218 1198
rect 3204 1041 3800 1155
rect 3204 1012 3218 1041
rect 2865 982 3218 1012
rect 2942 893 14872 933
rect 2942 888 13852 893
rect 2942 882 10413 888
rect 2942 860 7162 882
rect 664 838 7162 860
rect 664 474 696 838
rect 1202 504 7162 838
rect 7749 510 10413 882
rect 11000 515 13852 888
rect 14439 515 14872 893
rect 11000 510 14872 515
rect 7749 504 14872 510
rect 1202 474 14872 504
rect 664 456 14872 474
<< via1 >>
rect 2263 10817 2775 11264
rect 14397 10841 14842 11512
rect 1373 10489 1642 10646
rect 3320 10009 3623 10327
rect 1368 9726 1659 9848
rect 1808 9179 2110 9236
rect 704 8867 1200 9127
rect 1368 8099 1650 8304
rect 708 7300 1199 7565
rect 1808 7170 2108 7244
rect 1364 6565 1660 6697
rect 1378 5904 1635 6116
rect 2309 6126 2715 6454
rect 7191 5555 7795 6136
rect 10413 5589 11027 6136
rect 13849 5575 14463 6122
rect 3443 3979 3643 4179
rect 738 2141 1127 2862
rect 2877 1012 3204 1198
rect 696 474 1202 838
rect 7162 504 7749 882
rect 10413 510 11000 888
rect 13852 515 14439 893
<< metal2 >>
rect 2239 11264 2793 11285
rect 2239 10817 2263 11264
rect 2775 10817 2793 11264
rect 2239 10797 2793 10817
rect 1350 10646 1667 10669
rect 1350 10489 1373 10646
rect 1642 10489 1667 10646
rect 1350 10454 1667 10489
rect 6621 10379 6821 11552
rect 14370 11512 14880 11548
rect 14370 10841 14397 11512
rect 14842 10841 14880 11512
rect 14370 10809 14880 10841
rect 680 10327 3648 10343
rect 680 10109 3320 10327
rect 680 10026 706 10109
rect 1186 10026 3320 10109
rect 680 10009 3320 10026
rect 3623 10009 3648 10327
rect 680 9992 3648 10009
rect 1350 9886 1673 9903
rect 1350 9679 1368 9886
rect 1659 9679 1673 9886
rect 1350 9662 1673 9679
rect 1800 9314 2119 9324
rect 1800 9236 1809 9314
rect 1800 9179 1808 9236
rect 2111 9192 2119 9314
rect 2110 9179 2119 9192
rect 678 9127 1225 9151
rect 678 8867 704 9127
rect 1200 8867 1225 9127
rect 678 8842 1225 8867
rect 1353 8332 1669 8345
rect 1353 8099 1368 8332
rect 1650 8099 1669 8332
rect 1353 8074 1669 8099
rect 685 7565 1226 7595
rect 685 7300 708 7565
rect 1199 7300 1226 7565
rect 685 7276 1226 7300
rect 1800 7244 2119 7245
rect 1800 7049 1808 7244
rect 2108 7170 2119 7244
rect 2107 7049 2119 7170
rect 1800 7039 2119 7049
rect 3135 6764 3139 6809
rect 1350 6733 1667 6745
rect 1350 6697 1365 6733
rect 1655 6697 1667 6733
rect 1350 6565 1364 6697
rect 1660 6565 1667 6697
rect 1350 6537 1365 6565
rect 1655 6537 1667 6565
rect 3191 6564 5171 6609
rect 1350 6520 1667 6537
rect 2264 6455 2759 6496
rect 5464 6455 5982 6649
rect 2264 6454 5982 6455
rect 1351 6116 1668 6154
rect 1351 5904 1378 6116
rect 1635 5904 1668 6116
rect 2264 6126 2309 6454
rect 2715 6126 5982 6454
rect 2264 5992 2312 6126
rect 2712 5992 5982 6126
rect 2264 5937 5982 5992
rect 1351 5877 1668 5904
rect 1944 5770 3124 5899
rect 6703 5770 6903 6569
rect 1944 5759 6903 5770
rect 1944 5717 3376 5759
rect 1944 5304 2129 5717
rect 2906 5598 3376 5717
rect 3739 5598 6903 5759
rect 2906 5585 6903 5598
rect 7149 6195 7637 6625
rect 7149 6136 7834 6195
rect 7149 5555 7191 6136
rect 7795 5555 7834 6136
rect 10378 6187 10828 6655
rect 10378 6136 11063 6187
rect 14099 6174 14501 6640
rect 10378 5589 10413 6136
rect 11027 5589 11063 6136
rect 10378 5557 11063 5589
rect 13816 6122 14501 6174
rect 13816 5575 13849 6122
rect 14463 5575 14501 6122
rect 7149 5527 7834 5555
rect 13816 5542 14501 5575
rect 704 2862 1160 2891
rect 704 2141 738 2862
rect 1127 2141 1160 2862
rect 3045 2188 3089 5287
rect 704 2099 1160 2141
rect 3140 1307 3190 5437
rect 3443 5276 5433 5476
rect 3443 4179 3643 5276
rect 5233 5109 5433 5276
rect 3443 3970 3643 3979
rect 3140 1257 5167 1307
rect 2865 1198 3218 1217
rect 2865 1012 2877 1198
rect 3204 1012 3218 1198
rect 2865 997 3218 1012
rect 5465 957 5983 1368
rect 675 926 1224 952
rect 675 474 696 926
rect 1202 474 1224 926
rect 2724 852 5983 957
rect 675 452 1224 474
rect 2221 811 5983 852
rect 2221 468 2264 811
rect 2772 468 5983 811
rect 2221 439 5983 468
rect 6704 422 6904 1304
rect 7113 957 7600 1370
rect 7113 882 7798 957
rect 10519 949 10906 1412
rect 14100 966 14484 1373
rect 7113 504 7162 882
rect 7749 504 7798 882
rect 7113 457 7798 504
rect 10359 888 11044 949
rect 10359 510 10413 888
rect 11000 510 11044 888
rect 10359 460 11044 510
rect 13799 893 14484 966
rect 13799 515 13852 893
rect 14439 515 14484 893
rect 13799 460 14484 515
<< via2 >>
rect 2263 10817 2775 11264
rect 1373 10489 1642 10646
rect 14397 10841 14842 11512
rect 706 10026 1186 10109
rect 1368 9848 1659 9886
rect 1368 9726 1659 9848
rect 1368 9679 1659 9726
rect 1809 9236 2111 9314
rect 1809 9192 2110 9236
rect 2110 9192 2111 9236
rect 704 8867 1200 9127
rect 1368 8304 1650 8332
rect 1368 8099 1650 8304
rect 708 7300 1199 7565
rect 1808 7170 2107 7233
rect 1808 7049 2107 7170
rect 1365 6697 1655 6733
rect 1365 6565 1655 6697
rect 1365 6537 1655 6565
rect 1378 5904 1635 6116
rect 2312 6126 2712 6443
rect 2312 5992 2712 6126
rect 3376 5598 3739 5759
rect 738 2141 1127 2862
rect 2877 1012 3204 1198
rect 696 838 1202 926
rect 696 474 1202 838
rect 2264 468 2772 811
<< metal3 >>
rect 670 11349 1231 11558
rect 1350 11349 1670 11557
rect 1800 11553 2119 11556
rect 1800 11351 2120 11553
rect 675 10109 1229 11349
rect 675 10026 706 10109
rect 1186 10026 1229 10109
rect 675 9127 1229 10026
rect 675 8867 704 9127
rect 1200 8867 1229 9127
rect 675 7565 1229 8867
rect 675 7300 708 7565
rect 1199 7300 1229 7565
rect 675 2862 1229 7300
rect 675 2141 738 2862
rect 1127 2141 1229 2862
rect 675 1592 1229 2141
rect 1350 10646 1669 11349
rect 1350 10489 1373 10646
rect 1642 10489 1669 10646
rect 1350 9886 1669 10489
rect 1350 9679 1368 9886
rect 1659 9679 1669 9886
rect 1350 8332 1669 9679
rect 1350 8099 1368 8332
rect 1650 8099 1669 8332
rect 1350 6733 1669 8099
rect 1350 6537 1365 6733
rect 1655 6537 1669 6733
rect 1800 9314 2119 11351
rect 1800 9192 1809 9314
rect 2111 9192 2119 9314
rect 1800 7233 2119 9192
rect 1800 7049 1808 7233
rect 2107 7049 2119 7233
rect 1800 6648 2119 7049
rect 2239 11264 2793 11556
rect 2239 10817 2263 11264
rect 2775 10817 2793 11264
rect 1350 6116 1669 6537
rect 2239 6518 2793 10817
rect 14370 11512 14880 11548
rect 14370 10841 14397 11512
rect 14842 10841 14880 11512
rect 14370 10809 14880 10841
rect 1350 5904 1378 6116
rect 1635 5904 1669 6116
rect 2229 6443 2793 6518
rect 2229 5992 2312 6443
rect 2712 5992 2793 6443
rect 2229 5924 2793 5992
rect 675 926 1224 1592
rect 1350 1246 1669 5904
rect 1350 977 1377 1246
rect 1638 977 1669 1246
rect 1350 954 1669 977
rect 675 474 696 926
rect 1202 474 1224 926
rect 675 452 1224 474
rect 2239 811 2793 5924
rect 3358 5778 3753 5797
rect 3358 5545 3375 5778
rect 3733 5759 3753 5778
rect 3739 5598 3753 5759
rect 3733 5545 3753 5598
rect 3358 5528 3753 5545
rect 2865 1198 3218 1217
rect 2865 1012 2877 1198
rect 3204 1012 3218 1198
rect 2865 982 3218 1012
rect 2239 468 2264 811
rect 2772 468 2793 811
rect 2239 439 2793 468
<< via3 >>
rect 14397 10841 14842 11512
rect 1377 977 1638 1246
rect 3375 5759 3733 5778
rect 3375 5598 3376 5759
rect 3376 5598 3733 5759
rect 3375 5545 3733 5598
rect 2877 1012 3204 1198
<< metal4 >>
rect 14370 11512 14880 11548
rect 14370 10841 14397 11512
rect 14842 10841 14880 11512
rect 14370 10809 14880 10841
rect 3350 5849 3765 5879
rect 3350 5516 3375 5849
rect 3351 4956 3375 5516
rect 3733 4956 3765 5849
rect 3351 4927 3765 4956
rect 1350 1246 3220 1273
rect 1350 977 1377 1246
rect 1638 1198 3220 1246
rect 1638 1012 2877 1198
rect 3204 1012 3220 1198
rect 1638 977 3220 1012
rect 1350 954 3220 977
<< via4 >>
rect 3375 5778 3733 5849
rect 3375 5545 3733 5778
rect 3375 4956 3733 5545
<< metal5 >>
rect 3350 5849 3765 5879
rect 3350 5516 3375 5849
rect 3351 4956 3375 5516
rect 3733 4956 3765 5849
rect 3351 4927 3765 4956
use amp_via_4cut  amp_via_4cut_0
timestamp 1718240546
transform 0 1 11062 -1 0 21439
box 15948 -7932 16222 -7868
use amp_via_4cut  amp_via_4cut_1
timestamp 1718240546
transform 0 1 11065 -1 0 22776
box 15948 -7932 16222 -7868
use amp_via_4cut  amp_via_4cut_2
timestamp 1718240546
transform 0 1 10962 -1 0 21439
box 15948 -7932 16222 -7868
use amp_via_4cut  amp_via_4cut_3
timestamp 1718240546
transform 0 1 10967 -1 0 18142
box 15948 -7932 16222 -7868
use hold_cap_array  hold_cap_array_0
timestamp 1718240546
transform 0 1 29911 -1 0 13478
box 1925 -26553 13175 -15183
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_0 paramcells
timestamp 1718240546
transform 1 0 1386 0 1 6283
box -198 -198 198 198
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_1
timestamp 1718240546
transform 1 0 1351 0 1 10311
box -198 -198 198 198
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 875 0 -1 9840
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_1
timestamp 1715205430
transform 1 0 875 0 1 6584
box -66 -43 2178 1671
use balanced_switch  x1
timestamp 1718242347
transform -1 0 3080 0 -1 2783
box 301 -3111 2543 2130
use follower_amp  x2
timestamp 1718240546
transform 0 1 3724 1 0 1046
box 0 0 4377 11129
use follower_amp  x3
timestamp 1718240546
transform 0 1 3723 1 0 6294
box 0 0 4377 11129
<< labels >>
flabel metal2 6704 422 6904 622 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal3 2240 11349 2792 11556 0 FreeSans 1600 90 0 0 vss
port 5 nsew
flabel metal3 1800 11351 2120 11553 0 FreeSans 1600 90 0 0 dvdd
port 6 nsew
flabel metal3 1350 11349 1670 11557 0 FreeSans 1600 90 0 0 dvss
port 7 nsew
flabel metal3 670 11349 1231 11558 0 FreeSans 1600 90 0 0 vdd
port 2 nsew
flabel metal1 589 9358 786 9558 0 FreeSans 320 0 0 0 ena
port 8 nsew
flabel metal1 589 6842 789 7042 0 FreeSans 256 0 0 0 hold
port 3 nsew
flabel metal2 6621 11352 6821 11552 0 FreeSans 256 270 0 0 out
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 19469 11297
<< end >>
